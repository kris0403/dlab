`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:02:14 01/09/2016 
// Design Name: 
// Module Name:    rabiitgraph 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tuzki(
    input clk,
	 input[10:0] x,
	 input[10:0] y,
	 output reg word
    );
 wire [79:0] a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31,a32,a33,a34,a35,a36,a37,a38,a39,a40,a41,a42,a43,a44,a45,a46,a47,a48,a49,a50,a51,a52,a53,a54,a55,a56,a57,a58,a59,a60,a61,a62,a63,a64,a65,a66,a67,a68,a69,a70,a71,a72,a73,a74,a75,a76,a77,a78,a79,a80,a81,a82,a83,a84,a85,a86,a87,a88,a89,a90,a91,a92,a93,a94,a95,a96,a97,a98,a99,a100;



	assign a1  = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111;
	assign a2  = 80'b1000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000001;
	assign a3  = 80'b1000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000001;
	assign a4  = 80'b1000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000001;
	assign a5  = 80'b1000000000_0000000001_1111111111_0000000000_0000000001_1111111111_1000000000_0000000001;
	assign a6  = 80'b1000000000_0000000011_1111111111_1000000000_0000000001_1111111111_1000000000_0000000001;
	assign a7  = 80'b1000000000_0000000011_0000000001_1000000000_0000000011_0000000000_1100000000_0000000001;
	assign a8  = 80'b1000000000_0000000011_0000000000_1000000000_0000000011_0000000000_1100000000_0000000001;
	assign a9  = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a10 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a11 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a12 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a13 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a14 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a15 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a16 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a17 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a18 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a19 = 80'b1000000000_0000000011_0000000000_1100000000_0000000011_0000000000_1100000000_0000000001;
	assign a20 = 80'b1000000000_0000000011_1111111111_1111111111_1111111111_1111111111_1100000000_0000000001;
	assign a21 = 80'b1000000000_0000000111_1111111111_1111111111_1111111111_1111111111_1100000000_0000000001;
	assign a22 = 80'b1000000000_0000111100_0000000000_0000000000_0000000000_0000000011_1100000000_0000000001;
	assign a23 = 80'b1000000000_0001100000_0000000000_0000000000_0000000000_0000000011_1100000000_0000000001;
	assign a24 = 80'b1000000000_0011000000_0000000000_0000000000_0000000000_0000000000_1110000000_0000000001;
	assign a25 = 80'b1000000000_0110000000_0000000000_0000000000_0000000000_0000000000_0111000000_0000000001;
	assign a26 = 80'b1000000000_1100000000_0000000000_0000000000_0000000000_0000000000_0011000000_0000000001;
	assign a27 = 80'b1000000001_1000000000_0000000000_0000000000_0000000000_0000000000_0001100000_0000000001;
	assign a28 = 80'b1000000011_0000000000_0000000000_0000000000_0000000000_0000000000_0000110000_0000000001;
	assign a29 = 80'b1000000110_0000000000_0000000000_0000000000_0000000000_0000000000_0000110000_0000000001;
	assign a30 = 80'b1000001100_0000000000_0000000000_0000000000_0000000000_0000000000_0000011000_0000000001;
	assign a31 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a32 = 80'b1000111000_0011111111_1111111111_0000000000_1111111111_1111111111_0000001110_0000000001;
	assign a33 = 80'b1000111000_0011111111_1111111111_0000000000_1111111111_1111111111_0000001110_0000000001;
	assign a34 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a35 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a36 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a37 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a38 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a39 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a40 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a41 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a42 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a43 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a44 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a45 = 80'b1000111000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a46 = 80'b1000011000_0000000000_0000000000_0000000000_0000000000_0000000000_0000001110_0000000001;
	assign a47 = 80'b1000001100_0000000000_0000000000_0000000000_0000000000_0000000000_0000011100_0000000001;
	assign a48 = 80'b1000001100_0000000000_0000000000_0000000000_0000000000_0000000000_0000011000_0000000001;
	assign a49 = 80'b1000000110_0000000000_0000000000_0000000000_0000000000_0000000000_0000110000_0000000001;
	assign a50 = 80'b1000000011_0000000000_0000000000_0000000000_0000000000_0000000000_0001100000_0000000001;
	assign a51 = 80'b1000000001_1000000000_0000000000_0000000000_0000000000_0000000000_0011000000_0000000001;
	assign a52 = 80'b1000000000_1100000000_0000000000_0000000000_0000000000_0000000000_0110000000_0000000001;
	assign a53 = 80'b1000000000_0110000000_0000000000_0000000000_0000000000_0000000001_1000000000_0000000001;
	assign a54 = 80'b1000000000_0011111111_1111111111_0000000000_1111111111_1111111110_0000000000_0000000001;
	assign a55 = 80'b1000000000_0011111111_1111111111_0000000000_1111111111_1111111100_0000000000_0000000001;
	assign a56 = 80'b1000000000_1110000000_0000000000_0000000000_0000000000_0000000111_0000000000_0000000001;
	assign a57 = 80'b1000000001_1100000000_0000000000_0000000000_0000000000_0000000011_1000000000_0000000001;
	assign a58 = 80'b1000000011_1000000000_0000000000_0000000000_0000000000_0000000001_1100000000_0000000001;
	assign a59 = 80'b1000000111_0000000000_0000000000_0000000000_0000000000_0000000000_1110000000_0000000001;
	assign a60 = 80'b1000001110_0000001111_0000000000_0000000000_0000000000_1111000000_0111000000_0000000001;
	assign a61 = 80'b1000011100_0000001111_0000000000_0000000000_0000000000_1111000000_0011100000_0000000001;
	assign a62 = 80'b1000111000_0000011110_0000000000_0000000000_0000000000_0111000000_0001110000_0000000001;
	assign a63 = 80'b1000111000_0000011100_0000000000_0000000000_0000000000_0111000000_0001110000_0000000001;
	assign a64 = 80'b1000111000_0000011100_0000000000_0000000000_0000000000_0111000000_0001110000_0000000001;
	assign a65 = 80'b1000111000_0000011100_0000000000_0000000000_0000000000_0111000000_0001110000_0000000001;
	assign a66 = 80'b1000111000_0000111100_0000000000_0000000000_0000000000_1111000000_0001110000_0000000001;
	assign a67 = 80'b1000111000_0000111011_0000000000_0000000000_0000000011_0111000000_0001110000_0000000001;
	assign a68 = 80'b1000111000_0000111011_0000000000_0000000000_0000000011_0111000000_0001110000_0000000001;
	assign a69 = 80'b1000111000_0000111011_0000000000_0000000000_0000000011_0111000000_0001110000_0000000001;
	assign a70 = 80'b1000111000_0000111011_0000000000_0000000000_0000000011_0111000000_1111100000_0000000001;
	assign a71 = 80'b1000011111_1111111011_0000000000_0000000000_0000000011_0111111111_1111000000_0000000001;
	assign a72 = 80'b1000001111_1111100011_0000000000_0000000000_0000000011_0111111110_0000000000_0000000001;
	assign a73 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a74 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a75 = 80'b1000000000_0000000011_0000000000_0001001000_0000000011_0000000000_0000000000_0000000001;
	assign a76 = 80'b1000000000_0000000011_0000000000_0000110000_0000000011_0000000000_0000000000_0000000001;
	assign a77 = 80'b1000000000_0000000011_0000000000_0001001000_0000000011_0000000000_0000000000_0000000001;
	assign a78 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a79 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a80 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a81 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;	
	assign a82 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a83 = 80'b1000000000_0000000011_0000000000_0000000000_0000000011_0000000000_0000000000_0000000001;
	assign a84 = 80'b1000000000_0000000011_0000000011_0111111111_1100000011_0000000000_0000000000_0000000001;
	assign a85 = 80'b1000000000_0000000011_0000000011_0000000000_1100000011_0000000000_0000000000_0000000001;
	assign a86 = 80'b1000000000_0000000110_0000000011_0000000000_1100000001_1000000000_0000000000_0000000001;
	assign a87 = 80'b1000000000_0000000110_0000000011_0000000000_1100000001_1000000000_0000000000_0000000001;
	assign a88 = 80'b1000000000_0000001100_0000000011_0000000000_1100000000_1100000000_0000000000_0000000001;
	assign a89 = 80'b0000000000_0000011000_0000000011_0000000000_1100000000_0110000000_0000000000_0000000001;
	assign a90 = 80'b1000000000_0000110000_0000000011_0000000000_1100000000_0011000000_0000000000_0000000001;
	assign a91 = 80'b1000000000_0001100000_0000000011_0000000000_1100000000_0001100000_0000000000_0000000001;
	assign a92 = 80'b1000000000_0011000000_0000000011_0000000000_1100000000_0000110000_0000000000_0000000001;
	assign a93 = 80'b1000000000_0110000000_0000000011_0000000000_1100000000_0000011000_0000000000_0000000001;
	assign a94 = 80'b1000000000_0111111111_1111111111_0000000000_1111111111_1111101000_0000000000_0000000001;
	assign a95 = 80'b1111000011_1110000111_1111111111_1111111111_1111111111_1111111111_1111000011_1110000111;
	assign a96 = 80'b1111000011_1110000111_1111111111_1111111111_1111111111_1111111111_1111000011_1110000111;
	assign a97 = 80'b1000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000001;
	assign a98 = 80'b1000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000001;
	assign a99 = 80'b1000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000000_0000000001;
   assign a100 = 80'b1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111_1111111111;

always @(posedge clk)begin
	if(y >= 40 && y <= 140)begin
		case(y)
			40:begin
				case(x)
					290:word <= a1[0];
					289:word <= a1[1];
					287:word <= a1[2];
					286:word <= a1[3];
					285:word <= a1[4];
					284:word <= a1[5];
					283:word <= a1[6];
					282:word <= a1[7];
					281:word <= a1[8];
					280:word <= a1[9];
					279:word <= a1[10];
					278:word <= a1[11];
					277:word <= a1[12];
					276:word <= a1[13];
					275:word <= a1[14];
					274:word <= a1[15];
					273:word <= a1[16];
					272:word <= a1[17];
					271:word <= a1[18];
					270:word <= a1[19];
					269:word <= a1[20];
					268:word <= a1[21];
					267:word <= a1[22];
					266:word <= a1[23];
					265:word <= a1[24];
					264:word <= a1[25];
					263:word <= a1[26];
					262:word <= a1[27];
					261:word <= a1[28];
					260:word <= a1[29];
					259:word <= a1[30];
					258:word <= a1[31];
					257:word <= a1[32];
					256:word <= a1[33];
					255:word <= a1[34];
					254:word <= a1[35];
					253:word <= a1[36];
					252:word <= a1[37];
					251:word <= a1[38];
					250:word <= a1[39];
					249:word <= a1[40];
					248:word <= a1[41];
					247:word <= a1[42];
					246:word <= a1[43];
					245:word <= a1[44];
					244:word <= a1[45];
					243:word <= a1[46];
					242:word <= a1[47];
					241:word <= a1[48];
					240:word <= a1[49];
					239:word <= a1[50];
					238:word <= a1[51];
					237:word <= a1[52];
					236:word <= a1[53];
					235:word <= a1[54];
					234:word <= a1[55];
					233:word <= a1[56];
					232:word <= a1[57];
					231:word <= a1[58];
					230:word <= a1[59];
					229:word <= a1[60];
					228:word <= a1[61];
					227:word <= a1[62];
					226:word <= a1[63];
					225:word <= a1[64];
					224:word <= a1[65];
					223:word <= a1[66];
					222:word <= a1[67];
					221:word <= a1[68];
					220:word <= a1[69];
					219:word <= a1[70];
					218:word <= a1[71];
					217:word <= a1[72];
					216:word <= a1[73];
					215:word <= a1[74];
					214:word <= a1[75];
					213:word <= a1[76];
					212:word <= a1[77];
					211:word <= a1[78];
					default:word <= a1[79];
					endcase
				end
				41:begin
				case(x-100)
					290:word <= a2[0];
					289:word <= a2[1];
					287:word <= a2[2];
					286:word <= a2[3];
					285:word <= a2[4];
					284:word <= a2[5];
					283:word <= a2[6];
					282:word <= a2[7];
					281:word <= a2[8];
					280:word <= a2[9];
					279:word <= a2[10];
					278:word <= a2[11];
					277:word <= a2[12];
					276:word <= a2[13];
					275:word <= a2[14];
					274:word <= a2[15];
					273:word <= a2[16];
					272:word <= a2[17];
					271:word <= a2[18];
					270:word <= a2[19];
					269:word <= a2[20];
					268:word <= a2[21];
					267:word <= a2[22];
					266:word <= a2[23];
					265:word <= a2[24];
					264:word <= a2[25];
					263:word <= a2[26];
					262:word <= a2[27];
					261:word <= a2[28];
					260:word <= a2[29];
					259:word <= a2[30];
					258:word <= a2[31];
					257:word <= a2[32];
					256:word <= a2[33];
					255:word <= a2[34];
					254:word <= a2[35];
					253:word <= a2[36];
					252:word <= a2[37];
					251:word <= a2[38];
					250:word <= a2[39];
					249:word <= a2[40];
					248:word <= a2[41];
					247:word <= a2[42];
					246:word <= a2[43];
					245:word <= a2[44];
					244:word <= a2[45];
					243:word <= a2[46];
					242:word <= a2[47];
					241:word <= a2[48];
					240:word <= a2[49];
					239:word <= a2[50];
					238:word <= a2[51];
					237:word <= a2[52];
					236:word <= a2[53];
					235:word <= a2[54];
					234:word <= a2[55];
					233:word <= a2[56];
					232:word <= a2[57];
					231:word <= a2[58];
					230:word <= a2[59];
					229:word <= a2[60];
					228:word <= a2[61];
					227:word <= a2[62];
					226:word <= a2[63];
					225:word <= a2[64];
					224:word <= a2[65];
					223:word <= a2[66];
					222:word <= a2[67];
					221:word <= a2[68];
					220:word <= a2[69];
					219:word <= a2[70];
					218:word <= a2[71];
					217:word <= a2[72];
					216:word <= a2[73];
					215:word <= a2[74];
					214:word <= a2[75];
					213:word <= a2[76];
					212:word <= a2[77];
					211:word <= a2[78];
					default:word <= a2[79];
					endcase
				end
				43:begin
				case(x)
					290:word <= a3[0];
					289:word <= a3[1];
					287:word <= a3[2];
					286:word <= a3[3];
					285:word <= a3[4];
					284:word <= a3[5];
					283:word <= a3[6];
					282:word <= a3[7];
					281:word <= a3[8];
					280:word <= a3[9];
					279:word <= a3[10];
					278:word <= a3[11];
					277:word <= a3[12];
					276:word <= a3[13];
					275:word <= a3[14];
					274:word <= a3[15];
					273:word <= a3[16];
					272:word <= a3[17];
					271:word <= a3[18];
					270:word <= a3[19];
					269:word <= a3[20];
					268:word <= a3[21];
					267:word <= a3[22];
					266:word <= a3[23];
					265:word <= a3[24];
					264:word <= a3[25];
					263:word <= a3[26];
					262:word <= a3[27];
					261:word <= a3[28];
					260:word <= a3[29];
					259:word <= a3[30];
					258:word <= a3[31];
					257:word <= a3[32];
					256:word <= a3[33];
					255:word <= a3[34];
					254:word <= a3[35];
					253:word <= a3[36];
					252:word <= a3[37];
					251:word <= a3[38];
					250:word <= a3[39];
					249:word <= a3[40];
					248:word <= a3[41];
					247:word <= a3[42];
					246:word <= a3[43];
					245:word <= a3[44];
					244:word <= a3[45];
					243:word <= a3[46];
					242:word <= a3[47];
					241:word <= a3[48];
					240:word <= a3[49];
					239:word <= a3[50];
					238:word <= a3[51];
					237:word <= a3[52];
					236:word <= a3[53];
					235:word <= a3[54];
					234:word <= a3[55];
					233:word <= a3[56];
					232:word <= a3[57];
					231:word <= a3[58];
					230:word <= a3[59];
					229:word <= a3[60];
					228:word <= a3[61];
					227:word <= a3[62];
					226:word <= a3[63];
					225:word <= a3[64];
					224:word <= a3[65];
					223:word <= a3[66];
					222:word <= a3[67];
					221:word <= a3[68];
					220:word <= a3[69];
					219:word <= a3[70];
					218:word <= a3[71];
					217:word <= a3[72];
					216:word <= a3[73];
					215:word <= a3[74];
					214:word <= a3[75];
					213:word <= a3[76];
					212:word <= a3[77];
					211:word <= a3[78];
					default:word <= a3[79];
					endcase
				end
				44:begin
				case(x)
					290:word <= a4[0];
					289:word <= a4[1];
					287:word <= a4[2];
					286:word <= a4[3];
					285:word <= a4[4];
					284:word <= a4[5];
					283:word <= a4[6];
					282:word <= a4[7];
					281:word <= a4[8];
					280:word <= a4[9];
					279:word <= a4[10];
					278:word <= a4[11];
					277:word <= a4[12];
					276:word <= a4[13];
					275:word <= a4[14];
					274:word <= a4[15];
					273:word <= a4[16];
					272:word <= a4[17];
					271:word <= a4[18];
					270:word <= a4[19];
					269:word <= a4[20];
					268:word <= a4[21];
					267:word <= a4[22];
					266:word <= a4[23];
					265:word <= a4[24];
					264:word <= a4[25];
					263:word <= a4[26];
					262:word <= a4[27];
					261:word <= a4[28];
					260:word <= a4[29];
					259:word <= a4[30];
					258:word <= a4[31];
					257:word <= a4[32];
					256:word <= a4[33];
					255:word <= a4[34];
					254:word <= a4[35];
					253:word <= a4[36];
					252:word <= a4[37];
					251:word <= a4[38];
					250:word <= a4[39];
					249:word <= a4[40];
					248:word <= a4[41];
					247:word <= a4[42];
					246:word <= a4[43];
					245:word <= a4[44];
					244:word <= a4[45];
					243:word <= a4[46];
					242:word <= a4[47];
					241:word <= a4[48];
					240:word <= a4[49];
					239:word <= a4[50];
					238:word <= a4[51];
					237:word <= a4[52];
					236:word <= a4[53];
					235:word <= a4[54];
					234:word <= a4[55];
					233:word <= a4[56];
					232:word <= a4[57];
					231:word <= a4[58];
					230:word <= a4[59];
					229:word <= a4[60];
					228:word <= a4[61];
					227:word <= a4[62];
					226:word <= a4[63];
					225:word <= a4[64];
					224:word <= a4[65];
					223:word <= a4[66];
					222:word <= a4[67];
					221:word <= a4[68];
					220:word <= a4[69];
					219:word <= a4[70];
					218:word <= a4[71];
					217:word <= a4[72];
					216:word <= a4[73];
					215:word <= a4[74];
					214:word <= a4[75];
					213:word <= a4[76];
					212:word <= a4[77];
					211:word <= a4[78];
					default:word <= a4[79];
					endcase
				end
				45:begin
				case(x)
					290:word <= a5[0];
					289:word <= a5[1];
					287:word <= a5[2];
					286:word <= a5[3];
					285:word <= a5[4];
					284:word <= a5[5];
					283:word <= a5[6];
					282:word <= a5[7];
					281:word <= a5[8];
					280:word <= a5[9];
					279:word <= a5[10];
					278:word <= a5[11];
					277:word <= a5[12];
					276:word <= a5[13];
					275:word <= a5[14];
					274:word <= a5[15];
					273:word <= a5[16];
					272:word <= a5[17];
					271:word <= a5[18];
					270:word <= a5[19];
					269:word <= a5[20];
					268:word <= a5[21];
					267:word <= a5[22];
					266:word <= a5[23];
					265:word <= a5[24];
					264:word <= a5[25];
					263:word <= a5[26];
					262:word <= a5[27];
					261:word <= a5[28];
					260:word <= a5[29];
					259:word <= a5[30];
					258:word <= a5[31];
					257:word <= a5[32];
					256:word <= a5[33];
					255:word <= a5[34];
					254:word <= a5[35];
					253:word <= a5[36];
					252:word <= a5[37];
					251:word <= a5[38];
					250:word <= a5[39];
					249:word <= a5[40];
					248:word <= a5[41];
					247:word <= a5[42];
					246:word <= a5[43];
					245:word <= a5[44];
					244:word <= a5[45];
					243:word <= a5[46];
					242:word <= a5[47];
					241:word <= a5[48];
					240:word <= a5[49];
					239:word <= a5[50];
					238:word <= a5[51];
					237:word <= a5[52];
					236:word <= a5[53];
					235:word <= a5[54];
					234:word <= a5[55];
					233:word <= a5[56];
					232:word <= a5[57];
					231:word <= a5[58];
					230:word <= a5[59];
					229:word <= a5[60];
					228:word <= a5[61];
					227:word <= a5[62];
					226:word <= a5[63];
					225:word <= a5[64];
					224:word <= a5[65];
					223:word <= a5[66];
					222:word <= a5[67];
					221:word <= a5[68];
					220:word <= a5[69];
					219:word <= a5[70];
					218:word <= a5[71];
					217:word <= a5[72];
					216:word <= a5[73];
					215:word <= a5[74];
					214:word <= a5[75];
					213:word <= a5[76];
					212:word <= a5[77];
					211:word <= a5[78];
					default:word <= a5[79];
					endcase
				end
				46:begin
				case(x)
					290:word <= a6[0];
					289:word <= a6[1];
					287:word <= a6[2];
					286:word <= a6[3];
					285:word <= a6[4];
					284:word <= a6[5];
					283:word <= a6[6];
					282:word <= a6[7];
					281:word <= a6[8];
					280:word <= a6[9];
					279:word <= a6[10];
					278:word <= a6[11];
					277:word <= a6[12];
					276:word <= a6[13];
					275:word <= a6[14];
					274:word <= a6[15];
					273:word <= a6[16];
					272:word <= a6[17];
					271:word <= a6[18];
					270:word <= a6[19];
					269:word <= a6[20];
					268:word <= a6[21];
					267:word <= a6[22];
					266:word <= a6[23];
					265:word <= a6[24];
					264:word <= a6[25];
					263:word <= a6[26];
					262:word <= a6[27];
					261:word <= a6[28];
					260:word <= a6[29];
					259:word <= a6[30];
					258:word <= a6[31];
					257:word <= a6[32];
					256:word <= a6[33];
					255:word <= a6[34];
					254:word <= a6[35];
					253:word <= a6[36];
					252:word <= a6[37];
					251:word <= a6[38];
					250:word <= a6[39];
					249:word <= a6[40];
					248:word <= a6[41];
					247:word <= a6[42];
					246:word <= a6[43];
					245:word <= a6[44];
					244:word <= a6[45];
					243:word <= a6[46];
					242:word <= a6[47];
					241:word <= a6[48];
					240:word <= a6[49];
					239:word <= a6[50];
					238:word <= a6[51];
					237:word <= a6[52];
					236:word <= a6[53];
					235:word <= a6[54];
					234:word <= a6[55];
					233:word <= a6[56];
					232:word <= a6[57];
					231:word <= a6[58];
					230:word <= a6[59];
					229:word <= a6[60];
					228:word <= a6[61];
					227:word <= a6[62];
					226:word <= a6[63];
					225:word <= a6[64];
					224:word <= a6[65];
					223:word <= a6[66];
					222:word <= a6[67];
					221:word <= a6[68];
					220:word <= a6[69];
					219:word <= a6[70];
					218:word <= a6[71];
					217:word <= a6[72];
					216:word <= a6[73];
					215:word <= a6[74];
					214:word <= a6[75];
					213:word <= a6[76];
					212:word <= a6[77];
					211:word <= a6[78];
					default:word <= a6[79];
					endcase
				end
				47:begin
				case(x)
					290:word <= a7[0];
					289:word <= a7[1];
					287:word <= a7[2];
					286:word <= a7[3];
					285:word <= a7[4];
					284:word <= a7[5];
					283:word <= a7[6];
					282:word <= a7[7];
					281:word <= a7[8];
					280:word <= a7[9];
					279:word <= a7[10];
					278:word <= a7[11];
					277:word <= a7[12];
					276:word <= a7[13];
					275:word <= a7[14];
					274:word <= a7[15];
					273:word <= a7[16];
					272:word <= a7[17];
					271:word <= a7[18];
					270:word <= a7[19];
					269:word <= a7[20];
					268:word <= a7[21];
					267:word <= a7[22];
					266:word <= a7[23];
					265:word <= a7[24];
					264:word <= a7[25];
					263:word <= a7[26];
					262:word <= a7[27];
					261:word <= a7[28];
					260:word <= a7[29];
					259:word <= a7[30];
					258:word <= a7[31];
					257:word <= a7[32];
					256:word <= a7[33];
					255:word <= a7[34];
					254:word <= a7[35];
					253:word <= a7[36];
					252:word <= a7[37];
					251:word <= a7[38];
					250:word <= a7[39];
					249:word <= a7[40];
					248:word <= a7[41];
					247:word <= a7[42];
					246:word <= a7[43];
					245:word <= a7[44];
					244:word <= a7[45];
					243:word <= a7[46];
					242:word <= a7[47];
					241:word <= a7[48];
					240:word <= a7[49];
					239:word <= a7[50];
					238:word <= a7[51];
					237:word <= a7[52];
					236:word <= a7[53];
					235:word <= a7[54];
					234:word <= a7[55];
					233:word <= a7[56];
					232:word <= a7[57];
					231:word <= a7[58];
					230:word <= a7[59];
					229:word <= a7[60];
					228:word <= a7[61];
					227:word <= a7[62];
					226:word <= a7[63];
					225:word <= a7[64];
					224:word <= a7[65];
					223:word <= a7[66];
					222:word <= a7[67];
					221:word <= a7[68];
					220:word <= a7[69];
					219:word <= a7[70];
					218:word <= a7[71];
					217:word <= a7[72];
					216:word <= a7[73];
					215:word <= a7[74];
					214:word <= a7[75];
					213:word <= a7[76];
					212:word <= a7[77];
					211:word <= a7[78];
					default:word <= a7[79];
					endcase
				end
				48:begin
				case(x)
					290:word <= a8[0];
					289:word <= a8[1];
					287:word <= a8[2];
					286:word <= a8[3];
					285:word <= a8[4];
					284:word <= a8[5];
					283:word <= a8[6];
					282:word <= a8[7];
					281:word <= a8[8];
					280:word <= a8[9];
					279:word <= a8[10];
					278:word <= a8[11];
					277:word <= a8[12];
					276:word <= a8[13];
					275:word <= a8[14];
					274:word <= a8[15];
					273:word <= a8[16];
					272:word <= a8[17];
					271:word <= a8[18];
					270:word <= a8[19];
					269:word <= a8[20];
					268:word <= a8[21];
					267:word <= a8[22];
					266:word <= a8[23];
					265:word <= a8[24];
					264:word <= a8[25];
					263:word <= a8[26];
					262:word <= a8[27];
					261:word <= a8[28];
					260:word <= a8[29];
					259:word <= a8[30];
					258:word <= a8[31];
					257:word <= a8[32];
					256:word <= a8[33];
					255:word <= a8[34];
					254:word <= a8[35];
					253:word <= a8[36];
					252:word <= a8[37];
					251:word <= a8[38];
					250:word <= a8[39];
					249:word <= a8[40];
					248:word <= a8[41];
					247:word <= a8[42];
					246:word <= a8[43];
					245:word <= a8[44];
					244:word <= a8[45];
					243:word <= a8[46];
					242:word <= a8[47];
					241:word <= a8[48];
					240:word <= a8[49];
					239:word <= a8[50];
					238:word <= a8[51];
					237:word <= a8[52];
					236:word <= a8[53];
					235:word <= a8[54];
					234:word <= a8[55];
					233:word <= a8[56];
					232:word <= a8[57];
					231:word <= a8[58];
					230:word <= a8[59];
					229:word <= a8[60];
					228:word <= a8[61];
					227:word <= a8[62];
					226:word <= a8[63];
					225:word <= a8[64];
					224:word <= a8[65];
					223:word <= a8[66];
					222:word <= a8[67];
					221:word <= a8[68];
					220:word <= a8[69];
					219:word <= a8[70];
					218:word <= a8[71];
					217:word <= a8[72];
					216:word <= a8[73];
					215:word <= a8[74];
					214:word <= a8[75];
					213:word <= a8[76];
					212:word <= a8[77];
					211:word <= a8[78];
					default:word <= a8[79];
					endcase
				end
				49:begin
				case(x)
					290:word <= a9[0];
					289:word <= a9[1];
					287:word <= a9[2];
					286:word <= a9[3];
					285:word <= a9[4];
					284:word <= a9[5];
					283:word <= a9[6];
					282:word <= a9[7];
					281:word <= a9[8];
					280:word <= a9[9];
					279:word <= a9[10];
					278:word <= a9[11];
					277:word <= a9[12];
					276:word <= a9[13];
					275:word <= a9[14];
					274:word <= a9[15];
					273:word <= a9[16];
					272:word <= a9[17];
					271:word <= a9[18];
					270:word <= a9[19];
					269:word <= a9[20];
					268:word <= a9[21];
					267:word <= a9[22];
					266:word <= a9[23];
					265:word <= a9[24];
					264:word <= a9[25];
					263:word <= a9[26];
					262:word <= a9[27];
					261:word <= a9[28];
					260:word <= a9[29];
					259:word <= a9[30];
					258:word <= a9[31];
					257:word <= a9[32];
					256:word <= a9[33];
					255:word <= a9[34];
					254:word <= a9[35];
					253:word <= a9[36];
					252:word <= a9[37];
					251:word <= a9[38];
					250:word <= a9[39];
					249:word <= a9[40];
					248:word <= a9[41];
					247:word <= a9[42];
					246:word <= a9[43];
					245:word <= a9[44];
					244:word <= a9[45];
					243:word <= a9[46];
					242:word <= a9[47];
					241:word <= a9[48];
					240:word <= a9[49];
					239:word <= a9[50];
					238:word <= a9[51];
					237:word <= a9[52];
					236:word <= a9[53];
					235:word <= a9[54];
					234:word <= a9[55];
					233:word <= a9[56];
					232:word <= a9[57];
					231:word <= a9[58];
					230:word <= a9[59];
					229:word <= a9[60];
					228:word <= a9[61];
					227:word <= a9[62];
					226:word <= a9[63];
					225:word <= a9[64];
					224:word <= a9[65];
					223:word <= a9[66];
					222:word <= a9[67];
					221:word <= a9[68];
					220:word <= a9[69];
					219:word <= a9[70];
					218:word <= a9[71];
					217:word <= a9[72];
					216:word <= a9[73];
					215:word <= a9[74];
					214:word <= a9[75];
					213:word <= a9[76];
					212:word <= a9[77];
					211:word <= a9[78];
					default:word <= a9[79];
					endcase
				end
				50:begin
				case(x)
					290:word <= a10[0];
					289:word <= a10[1];
					287:word <= a10[2];
					286:word <= a10[3];
					285:word <= a10[4];
					284:word <= a10[5];
					283:word <= a10[6];
					282:word <= a10[7];
					281:word <= a10[8];
					280:word <= a10[9];
					279:word <= a10[10];
					278:word <= a10[11];
					277:word <= a10[12];
					276:word <= a10[13];
					275:word <= a10[14];
					274:word <= a10[15];
					273:word <= a10[16];
					272:word <= a10[17];
					271:word <= a10[18];
					270:word <= a10[19];
					269:word <= a10[20];
					268:word <= a10[21];
					267:word <= a10[22];
					266:word <= a10[23];
					265:word <= a10[24];
					264:word <= a10[25];
					263:word <= a10[26];
					262:word <= a10[27];
					261:word <= a10[28];
					260:word <= a10[29];
					259:word <= a10[30];
					258:word <= a10[31];
					257:word <= a10[32];
					256:word <= a10[33];
					255:word <= a10[34];
					254:word <= a10[35];
					253:word <= a10[36];
					252:word <= a10[37];
					251:word <= a10[38];
					250:word <= a10[39];
					249:word <= a10[40];
					248:word <= a10[41];
					247:word <= a10[42];
					246:word <= a10[43];
					245:word <= a10[44];
					244:word <= a10[45];
					243:word <= a10[46];
					242:word <= a10[47];
					241:word <= a10[48];
					240:word <= a10[49];
					239:word <= a10[50];
					238:word <= a10[51];
					237:word <= a10[52];
					236:word <= a10[53];
					235:word <= a10[54];
					234:word <= a10[55];
					233:word <= a10[56];
					232:word <= a10[57];
					231:word <= a10[58];
					230:word <= a10[59];
					229:word <= a10[60];
					228:word <= a10[61];
					227:word <= a10[62];
					226:word <= a10[63];
					225:word <= a10[64];
					224:word <= a10[65];
					223:word <= a10[66];
					222:word <= a10[67];
					221:word <= a10[68];
					220:word <= a10[69];
					219:word <= a10[70];
					218:word <= a10[71];
					217:word <= a10[72];
					216:word <= a10[73];
					215:word <= a10[74];
					214:word <= a10[75];
					213:word <= a10[76];
					212:word <= a10[77];
					211:word <= a10[78];
					default:word <= a10[79];
					endcase
				end
				51:begin
				case(x)
					290:word <= a11[0];
					289:word <= a11[1];
					287:word <= a11[2];
					286:word <= a11[3];
					285:word <= a11[4];
					284:word <= a11[5];
					283:word <= a11[6];
					282:word <= a11[7];
					281:word <= a11[8];
					280:word <= a11[9];
					279:word <= a11[10];
					278:word <= a11[11];
					277:word <= a11[12];
					276:word <= a11[13];
					275:word <= a11[14];
					274:word <= a11[15];
					273:word <= a11[16];
					272:word <= a11[17];
					271:word <= a11[18];
					270:word <= a11[19];
					269:word <= a11[20];
					268:word <= a11[21];
					267:word <= a11[22];
					266:word <= a11[23];
					265:word <= a11[24];
					264:word <= a11[25];
					263:word <= a11[26];
					262:word <= a11[27];
					261:word <= a11[28];
					260:word <= a11[29];
					259:word <= a11[30];
					258:word <= a11[31];
					257:word <= a11[32];
					256:word <= a11[33];
					255:word <= a11[34];
					254:word <= a11[35];
					253:word <= a11[36];
					252:word <= a11[37];
					251:word <= a11[38];
					250:word <= a11[39];
					249:word <= a11[40];
					248:word <= a11[41];
					247:word <= a11[42];
					246:word <= a11[43];
					245:word <= a11[44];
					244:word <= a11[45];
					243:word <= a11[46];
					242:word <= a11[47];
					241:word <= a11[48];
					240:word <= a11[49];
					239:word <= a11[50];
					238:word <= a11[51];
					237:word <= a11[52];
					236:word <= a11[53];
					235:word <= a11[54];
					234:word <= a11[55];
					233:word <= a11[56];
					232:word <= a11[57];
					231:word <= a11[58];
					230:word <= a11[59];
					229:word <= a11[60];
					228:word <= a11[61];
					227:word <= a11[62];
					226:word <= a11[63];
					225:word <= a11[64];
					224:word <= a11[65];
					223:word <= a11[66];
					222:word <= a11[67];
					221:word <= a11[68];
					220:word <= a11[69];
					219:word <= a11[70];
					218:word <= a11[71];
					217:word <= a11[72];
					216:word <= a11[73];
					215:word <= a11[74];
					214:word <= a11[75];
					213:word <= a11[76];
					212:word <= a11[77];
					211:word <= a11[78];
					default:word <= a11[79];
					endcase
				end
				52:begin
				case(x)
					290:word <= a12[0];
					289:word <= a12[1];
					287:word <= a12[2];
					286:word <= a12[3];
					285:word <= a12[4];
					284:word <= a12[5];
					283:word <= a12[6];
					282:word <= a12[7];
					281:word <= a12[8];
					280:word <= a12[9];
					279:word <= a12[10];
					278:word <= a12[11];
					277:word <= a12[12];
					276:word <= a12[13];
					275:word <= a12[14];
					274:word <= a12[15];
					273:word <= a12[16];
					272:word <= a12[17];
					271:word <= a12[18];
					270:word <= a12[19];
					269:word <= a12[20];
					268:word <= a12[21];
					267:word <= a12[22];
					266:word <= a12[23];
					265:word <= a12[24];
					264:word <= a12[25];
					263:word <= a12[26];
					262:word <= a12[27];
					261:word <= a12[28];
					260:word <= a12[29];
					259:word <= a12[30];
					258:word <= a12[31];
					257:word <= a12[32];
					256:word <= a12[33];
					255:word <= a12[34];
					254:word <= a12[35];
					253:word <= a12[36];
					252:word <= a12[37];
					251:word <= a12[38];
					250:word <= a12[39];
					249:word <= a12[40];
					248:word <= a12[41];
					247:word <= a12[42];
					246:word <= a12[43];
					245:word <= a12[44];
					244:word <= a12[45];
					243:word <= a12[46];
					242:word <= a12[47];
					241:word <= a12[48];
					240:word <= a12[49];
					239:word <= a12[50];
					238:word <= a12[51];
					237:word <= a12[52];
					236:word <= a12[53];
					235:word <= a12[54];
					234:word <= a12[55];
					233:word <= a12[56];
					232:word <= a12[57];
					231:word <= a12[58];
					230:word <= a12[59];
					229:word <= a12[60];
					228:word <= a12[61];
					227:word <= a12[62];
					226:word <= a12[63];
					225:word <= a12[64];
					224:word <= a12[65];
					223:word <= a12[66];
					222:word <= a12[67];
					221:word <= a12[68];
					220:word <= a12[69];
					219:word <= a12[70];
					218:word <= a12[71];
					217:word <= a12[72];
					216:word <= a12[73];
					215:word <= a12[74];
					214:word <= a12[75];
					213:word <= a12[76];
					212:word <= a12[77];
					211:word <= a12[78];
					default:word <= a12[79];
					endcase
				end
				53:begin
				case(x)
					290:word <= a13[0];
					289:word <= a13[1];
					287:word <= a13[2];
					286:word <= a13[3];
					285:word <= a13[4];
					284:word <= a13[5];
					283:word <= a13[6];
					282:word <= a13[7];
					281:word <= a13[8];
					280:word <= a13[9];
					279:word <= a13[10];
					278:word <= a13[11];
					277:word <= a13[12];
					276:word <= a13[13];
					275:word <= a13[14];
					274:word <= a13[15];
					273:word <= a13[16];
					272:word <= a13[17];
					271:word <= a13[18];
					270:word <= a13[19];
					269:word <= a13[20];
					268:word <= a13[21];
					267:word <= a13[22];
					266:word <= a13[23];
					265:word <= a13[24];
					264:word <= a13[25];
					263:word <= a13[26];
					262:word <= a13[27];
					261:word <= a13[28];
					260:word <= a13[29];
					259:word <= a13[30];
					258:word <= a13[31];
					257:word <= a13[32];
					256:word <= a13[33];
					255:word <= a13[34];
					254:word <= a13[35];
					253:word <= a13[36];
					252:word <= a13[37];
					251:word <= a13[38];
					250:word <= a13[39];
					249:word <= a13[40];
					248:word <= a13[41];
					247:word <= a13[42];
					246:word <= a13[43];
					245:word <= a13[44];
					244:word <= a13[45];
					243:word <= a13[46];
					242:word <= a13[47];
					241:word <= a13[48];
					240:word <= a13[49];
					239:word <= a13[50];
					238:word <= a13[51];
					237:word <= a13[52];
					236:word <= a13[53];
					235:word <= a13[54];
					234:word <= a13[55];
					233:word <= a13[56];
					232:word <= a13[57];
					231:word <= a13[58];
					230:word <= a13[59];
					229:word <= a13[60];
					228:word <= a13[61];
					227:word <= a13[62];
					226:word <= a13[63];
					225:word <= a13[64];
					224:word <= a13[65];
					223:word <= a13[66];
					222:word <= a13[67];
					221:word <= a13[68];
					220:word <= a13[69];
					219:word <= a13[70];
					218:word <= a13[71];
					217:word <= a13[72];
					216:word <= a13[73];
					215:word <= a13[74];
					214:word <= a13[75];
					213:word <= a13[76];
					212:word <= a13[77];
					211:word <= a13[78];
					default:word <= a13[79];
					endcase
				end
				54:begin
				case(x)
					290:word <= a14[0];
					289:word <= a14[1];
					287:word <= a14[2];
					286:word <= a14[3];
					285:word <= a14[4];
					284:word <= a14[5];
					283:word <= a14[6];
					282:word <= a14[7];
					281:word <= a14[8];
					280:word <= a14[9];
					279:word <= a14[10];
					278:word <= a14[11];
					277:word <= a14[12];
					276:word <= a14[13];
					275:word <= a14[14];
					274:word <= a14[15];
					273:word <= a14[16];
					272:word <= a14[17];
					271:word <= a14[18];
					270:word <= a14[19];
					269:word <= a14[20];
					268:word <= a14[21];
					267:word <= a14[22];
					266:word <= a14[23];
					265:word <= a14[24];
					264:word <= a14[25];
					263:word <= a14[26];
					262:word <= a14[27];
					261:word <= a14[28];
					260:word <= a14[29];
					259:word <= a14[30];
					258:word <= a14[31];
					257:word <= a14[32];
					256:word <= a14[33];
					255:word <= a14[34];
					254:word <= a14[35];
					253:word <= a14[36];
					252:word <= a14[37];
					251:word <= a14[38];
					250:word <= a14[39];
					249:word <= a14[40];
					248:word <= a14[41];
					247:word <= a14[42];
					246:word <= a14[43];
					245:word <= a14[44];
					244:word <= a14[45];
					243:word <= a14[46];
					242:word <= a14[47];
					241:word <= a14[48];
					240:word <= a14[49];
					239:word <= a14[50];
					238:word <= a14[51];
					237:word <= a14[52];
					236:word <= a14[53];
					235:word <= a14[54];
					234:word <= a14[55];
					233:word <= a14[56];
					232:word <= a14[57];
					231:word <= a14[58];
					230:word <= a14[59];
					229:word <= a14[60];
					228:word <= a14[61];
					227:word <= a14[62];
					226:word <= a14[63];
					225:word <= a14[64];
					224:word <= a14[65];
					223:word <= a14[66];
					222:word <= a14[67];
					221:word <= a14[68];
					220:word <= a14[69];
					219:word <= a14[70];
					218:word <= a14[71];
					217:word <= a14[72];
					216:word <= a14[73];
					215:word <= a14[74];
					214:word <= a14[75];
					213:word <= a14[76];
					212:word <= a14[77];
					211:word <= a14[78];
					default:word <= a14[79];
					endcase
				end
				55:begin
				case(x)
					290:word <= a15[0];
					289:word <= a15[1];
					287:word <= a15[2];
					286:word <= a15[3];
					285:word <= a15[4];
					284:word <= a15[5];
					283:word <= a15[6];
					282:word <= a15[7];
					281:word <= a15[8];
					280:word <= a15[9];
					279:word <= a15[10];
					278:word <= a15[11];
					277:word <= a15[12];
					276:word <= a15[13];
					275:word <= a15[14];
					274:word <= a15[15];
					273:word <= a15[16];
					272:word <= a15[17];
					271:word <= a15[18];
					270:word <= a15[19];
					269:word <= a15[20];
					268:word <= a15[21];
					267:word <= a15[22];
					266:word <= a15[23];
					265:word <= a15[24];
					264:word <= a15[25];
					263:word <= a15[26];
					262:word <= a15[27];
					261:word <= a15[28];
					260:word <= a15[29];
					259:word <= a15[30];
					258:word <= a15[31];
					257:word <= a15[32];
					256:word <= a15[33];
					255:word <= a15[34];
					254:word <= a15[35];
					253:word <= a15[36];
					252:word <= a15[37];
					251:word <= a15[38];
					250:word <= a15[39];
					249:word <= a15[40];
					248:word <= a15[41];
					247:word <= a15[42];
					246:word <= a15[43];
					245:word <= a15[44];
					244:word <= a15[45];
					243:word <= a15[46];
					242:word <= a15[47];
					241:word <= a15[48];
					240:word <= a15[49];
					239:word <= a15[50];
					238:word <= a15[51];
					237:word <= a15[52];
					236:word <= a15[53];
					235:word <= a15[54];
					234:word <= a15[55];
					233:word <= a15[56];
					232:word <= a15[57];
					231:word <= a15[58];
					230:word <= a15[59];
					229:word <= a15[60];
					228:word <= a15[61];
					227:word <= a15[62];
					226:word <= a15[63];
					225:word <= a15[64];
					224:word <= a15[65];
					223:word <= a15[66];
					222:word <= a15[67];
					221:word <= a15[68];
					220:word <= a15[69];
					219:word <= a15[70];
					218:word <= a15[71];
					217:word <= a15[72];
					216:word <= a15[73];
					215:word <= a15[74];
					214:word <= a15[75];
					213:word <= a15[76];
					212:word <= a15[77];
					211:word <= a15[78];
					default:word <= a15[79];
					endcase
				end
				56:begin
				case(x)
					290:word <= a16[0];
					289:word <= a16[1];
					287:word <= a16[2];
					286:word <= a16[3];
					285:word <= a16[4];
					284:word <= a16[5];
					283:word <= a16[6];
					282:word <= a16[7];
					281:word <= a16[8];
					280:word <= a16[9];
					279:word <= a16[10];
					278:word <= a16[11];
					277:word <= a16[12];
					276:word <= a16[13];
					275:word <= a16[14];
					274:word <= a16[15];
					273:word <= a16[16];
					272:word <= a16[17];
					271:word <= a16[18];
					270:word <= a16[19];
					269:word <= a16[20];
					268:word <= a16[21];
					267:word <= a16[22];
					266:word <= a16[23];
					265:word <= a16[24];
					264:word <= a16[25];
					263:word <= a16[26];
					262:word <= a16[27];
					261:word <= a16[28];
					260:word <= a16[29];
					259:word <= a16[30];
					258:word <= a16[31];
					257:word <= a16[32];
					256:word <= a16[33];
					255:word <= a16[34];
					254:word <= a16[35];
					253:word <= a16[36];
					252:word <= a16[37];
					251:word <= a16[38];
					250:word <= a16[39];
					249:word <= a16[40];
					248:word <= a16[41];
					247:word <= a16[42];
					246:word <= a16[43];
					245:word <= a16[44];
					244:word <= a16[45];
					243:word <= a16[46];
					242:word <= a16[47];
					241:word <= a16[48];
					240:word <= a16[49];
					239:word <= a16[50];
					238:word <= a16[51];
					237:word <= a16[52];
					236:word <= a16[53];
					235:word <= a16[54];
					234:word <= a16[55];
					233:word <= a16[56];
					232:word <= a16[57];
					231:word <= a16[58];
					230:word <= a16[59];
					229:word <= a16[60];
					228:word <= a16[61];
					227:word <= a16[62];
					226:word <= a16[63];
					225:word <= a16[64];
					224:word <= a16[65];
					223:word <= a16[66];
					222:word <= a16[67];
					221:word <= a16[68];
					220:word <= a16[69];
					219:word <= a16[70];
					218:word <= a16[71];
					217:word <= a16[72];
					216:word <= a16[73];
					215:word <= a16[74];
					214:word <= a16[75];
					213:word <= a16[76];
					212:word <= a16[77];
					211:word <= a16[78];
					default:word <= a16[79];
					endcase
				end
				57:begin
				case(x)
					290:word <= a17[0];
					289:word <= a17[1];
					287:word <= a17[2];
					286:word <= a17[3];
					285:word <= a17[4];
					284:word <= a17[5];
					283:word <= a17[6];
					282:word <= a17[7];
					281:word <= a17[8];
					280:word <= a17[9];
					279:word <= a17[10];
					278:word <= a17[11];
					277:word <= a17[12];
					276:word <= a17[13];
					275:word <= a17[14];
					274:word <= a17[15];
					273:word <= a17[16];
					272:word <= a17[17];
					271:word <= a17[18];
					270:word <= a17[19];
					269:word <= a17[20];
					268:word <= a17[21];
					267:word <= a17[22];
					266:word <= a17[23];
					265:word <= a17[24];
					264:word <= a17[25];
					263:word <= a17[26];
					262:word <= a17[27];
					261:word <= a17[28];
					260:word <= a17[29];
					259:word <= a17[30];
					258:word <= a17[31];
					257:word <= a17[32];
					256:word <= a17[33];
					255:word <= a17[34];
					254:word <= a17[35];
					253:word <= a17[36];
					252:word <= a17[37];
					251:word <= a17[38];
					250:word <= a17[39];
					249:word <= a17[40];
					248:word <= a17[41];
					247:word <= a17[42];
					246:word <= a17[43];
					245:word <= a17[44];
					244:word <= a17[45];
					243:word <= a17[46];
					242:word <= a17[47];
					241:word <= a17[48];
					240:word <= a17[49];
					239:word <= a17[50];
					238:word <= a17[51];
					237:word <= a17[52];
					236:word <= a17[53];
					235:word <= a17[54];
					234:word <= a17[55];
					233:word <= a17[56];
					232:word <= a17[57];
					231:word <= a17[58];
					230:word <= a17[59];
					229:word <= a17[60];
					228:word <= a17[61];
					227:word <= a17[62];
					226:word <= a17[63];
					225:word <= a17[64];
					224:word <= a17[65];
					223:word <= a17[66];
					222:word <= a17[67];
					221:word <= a17[68];
					220:word <= a17[69];
					219:word <= a17[70];
					218:word <= a17[71];
					217:word <= a17[72];
					216:word <= a17[73];
					215:word <= a17[74];
					214:word <= a17[75];
					213:word <= a17[76];
					212:word <= a17[77];
					211:word <= a17[78];
					default:word <= a17[79];
					endcase
				end
				58:begin
				case(x)
					290:word <= a18[0];
					289:word <= a18[1];
					287:word <= a18[2];
					286:word <= a18[3];
					285:word <= a18[4];
					284:word <= a18[5];
					283:word <= a18[6];
					282:word <= a18[7];
					281:word <= a18[8];
					280:word <= a18[9];
					279:word <= a18[10];
					278:word <= a18[11];
					277:word <= a18[12];
					276:word <= a18[13];
					275:word <= a18[14];
					274:word <= a18[15];
					273:word <= a18[16];
					272:word <= a18[17];
					271:word <= a18[18];
					270:word <= a18[19];
					269:word <= a18[20];
					268:word <= a18[21];
					267:word <= a18[22];
					266:word <= a18[23];
					265:word <= a18[24];
					264:word <= a18[25];
					263:word <= a18[26];
					262:word <= a18[27];
					261:word <= a18[28];
					260:word <= a18[29];
					259:word <= a18[30];
					258:word <= a18[31];
					257:word <= a18[32];
					256:word <= a18[33];
					255:word <= a18[34];
					254:word <= a18[35];
					253:word <= a18[36];
					252:word <= a18[37];
					251:word <= a18[38];
					250:word <= a18[39];
					249:word <= a18[40];
					248:word <= a18[41];
					247:word <= a18[42];
					246:word <= a18[43];
					245:word <= a18[44];
					244:word <= a18[45];
					243:word <= a18[46];
					242:word <= a18[47];
					241:word <= a18[48];
					240:word <= a18[49];
					239:word <= a18[50];
					238:word <= a18[51];
					237:word <= a18[52];
					236:word <= a18[53];
					235:word <= a18[54];
					234:word <= a18[55];
					233:word <= a18[56];
					232:word <= a18[57];
					231:word <= a18[58];
					230:word <= a18[59];
					229:word <= a18[60];
					228:word <= a18[61];
					227:word <= a18[62];
					226:word <= a18[63];
					225:word <= a18[64];
					224:word <= a18[65];
					223:word <= a18[66];
					222:word <= a18[67];
					221:word <= a18[68];
					220:word <= a18[69];
					219:word <= a18[70];
					218:word <= a18[71];
					217:word <= a18[72];
					216:word <= a18[73];
					215:word <= a18[74];
					214:word <= a18[75];
					213:word <= a18[76];
					212:word <= a18[77];
					211:word <= a18[78];
					default:word <= a18[79];
					endcase
				end
				59:begin
				case(x)
					290:word <= a19[0];
					289:word <= a19[1];
					287:word <= a19[2];
					286:word <= a19[3];
					285:word <= a19[4];
					284:word <= a19[5];
					283:word <= a19[6];
					282:word <= a19[7];
					281:word <= a19[8];
					280:word <= a19[9];
					279:word <= a19[10];
					278:word <= a19[11];
					277:word <= a19[12];
					276:word <= a19[13];
					275:word <= a19[14];
					274:word <= a19[15];
					273:word <= a19[16];
					272:word <= a19[17];
					271:word <= a19[18];
					270:word <= a19[19];
					269:word <= a19[20];
					268:word <= a19[21];
					267:word <= a19[22];
					266:word <= a19[23];
					265:word <= a19[24];
					264:word <= a19[25];
					263:word <= a19[26];
					262:word <= a19[27];
					261:word <= a19[28];
					260:word <= a19[29];
					259:word <= a19[30];
					258:word <= a19[31];
					257:word <= a19[32];
					256:word <= a19[33];
					255:word <= a19[34];
					254:word <= a19[35];
					253:word <= a19[36];
					252:word <= a19[37];
					251:word <= a19[38];
					250:word <= a19[39];
					249:word <= a19[40];
					248:word <= a19[41];
					247:word <= a19[42];
					246:word <= a19[43];
					245:word <= a19[44];
					244:word <= a19[45];
					243:word <= a19[46];
					242:word <= a19[47];
					241:word <= a19[48];
					240:word <= a19[49];
					239:word <= a19[50];
					238:word <= a19[51];
					237:word <= a19[52];
					236:word <= a19[53];
					235:word <= a19[54];
					234:word <= a19[55];
					233:word <= a19[56];
					232:word <= a19[57];
					231:word <= a19[58];
					230:word <= a19[59];
					229:word <= a19[60];
					228:word <= a19[61];
					227:word <= a19[62];
					226:word <= a19[63];
					225:word <= a19[64];
					224:word <= a19[65];
					223:word <= a19[66];
					222:word <= a19[67];
					221:word <= a19[68];
					220:word <= a19[69];
					219:word <= a19[70];
					218:word <= a19[71];
					217:word <= a19[72];
					216:word <= a19[73];
					215:word <= a19[74];
					214:word <= a19[75];
					213:word <= a19[76];
					212:word <= a19[77];
					211:word <= a19[78];
					default:word <= a19[79];
					endcase
				end
				60:begin
				case(x)
					290:word <= a20[0];
					289:word <= a20[1];
					287:word <= a20[2];
					286:word <= a20[3];
					285:word <= a20[4];
					284:word <= a20[5];
					283:word <= a20[6];
					282:word <= a20[7];
					281:word <= a20[8];
					280:word <= a20[9];
					279:word <= a20[10];
					278:word <= a20[11];
					277:word <= a20[12];
					276:word <= a20[13];
					275:word <= a20[14];
					274:word <= a20[15];
					273:word <= a20[16];
					272:word <= a20[17];
					271:word <= a20[18];
					270:word <= a20[19];
					269:word <= a20[20];
					268:word <= a20[21];
					267:word <= a20[22];
					266:word <= a20[23];
					265:word <= a20[24];
					264:word <= a20[25];
					263:word <= a20[26];
					262:word <= a20[27];
					261:word <= a20[28];
					260:word <= a20[29];
					259:word <= a20[30];
					258:word <= a20[31];
					257:word <= a20[32];
					256:word <= a20[33];
					255:word <= a20[34];
					254:word <= a20[35];
					253:word <= a20[36];
					252:word <= a20[37];
					251:word <= a20[38];
					250:word <= a20[39];
					249:word <= a20[40];
					248:word <= a20[41];
					247:word <= a20[42];
					246:word <= a20[43];
					245:word <= a20[44];
					244:word <= a20[45];
					243:word <= a20[46];
					242:word <= a20[47];
					241:word <= a20[48];
					240:word <= a20[49];
					239:word <= a20[50];
					238:word <= a20[51];
					237:word <= a20[52];
					236:word <= a20[53];
					235:word <= a20[54];
					234:word <= a20[55];
					233:word <= a20[56];
					232:word <= a20[57];
					231:word <= a20[58];
					230:word <= a20[59];
					229:word <= a20[60];
					228:word <= a20[61];
					227:word <= a20[62];
					226:word <= a20[63];
					225:word <= a20[64];
					224:word <= a20[65];
					223:word <= a20[66];
					222:word <= a20[67];
					221:word <= a20[68];
					220:word <= a20[69];
					219:word <= a20[70];
					218:word <= a20[71];
					217:word <= a20[72];
					216:word <= a20[73];
					215:word <= a20[74];
					214:word <= a20[75];
					213:word <= a20[76];
					212:word <= a20[77];
					211:word <= a20[78];
					default:word <= a20[79];
					endcase
				end
				61:begin
				case(x)
					290:word <= a21[0];
					289:word <= a21[1];
					287:word <= a21[2];
					286:word <= a21[3];
					285:word <= a21[4];
					284:word <= a21[5];
					283:word <= a21[6];
					282:word <= a21[7];
					281:word <= a21[8];
					280:word <= a21[9];
					279:word <= a21[10];
					278:word <= a21[11];
					277:word <= a21[12];
					276:word <= a21[13];
					275:word <= a21[14];
					274:word <= a21[15];
					273:word <= a21[16];
					272:word <= a21[17];
					271:word <= a21[18];
					270:word <= a21[19];
					269:word <= a21[20];
					268:word <= a21[21];
					267:word <= a21[22];
					266:word <= a21[23];
					265:word <= a21[24];
					264:word <= a21[25];
					263:word <= a21[26];
					262:word <= a21[27];
					261:word <= a21[28];
					260:word <= a21[29];
					259:word <= a21[30];
					258:word <= a21[31];
					257:word <= a21[32];
					256:word <= a21[33];
					255:word <= a21[34];
					254:word <= a21[35];
					253:word <= a21[36];
					252:word <= a21[37];
					251:word <= a21[38];
					250:word <= a21[39];
					249:word <= a21[40];
					248:word <= a21[41];
					247:word <= a21[42];
					246:word <= a21[43];
					245:word <= a21[44];
					244:word <= a21[45];
					243:word <= a21[46];
					242:word <= a21[47];
					241:word <= a21[48];
					240:word <= a21[49];
					239:word <= a21[50];
					238:word <= a21[51];
					237:word <= a21[52];
					236:word <= a21[53];
					235:word <= a21[54];
					234:word <= a21[55];
					233:word <= a21[56];
					232:word <= a21[57];
					231:word <= a21[58];
					230:word <= a21[59];
					229:word <= a21[60];
					228:word <= a21[61];
					227:word <= a21[62];
					226:word <= a21[63];
					225:word <= a21[64];
					224:word <= a21[65];
					223:word <= a21[66];
					222:word <= a21[67];
					221:word <= a21[68];
					220:word <= a21[69];
					219:word <= a21[70];
					218:word <= a21[71];
					217:word <= a21[72];
					216:word <= a21[73];
					215:word <= a21[74];
					214:word <= a21[75];
					213:word <= a21[76];
					212:word <= a21[77];
					211:word <= a21[78];
					default:word <= a21[79];
					endcase
				end
				62:begin
				case(x)
					290:word <= a22[0];
					289:word <= a22[1];
					287:word <= a22[2];
					286:word <= a22[3];
					285:word <= a22[4];
					284:word <= a22[5];
					283:word <= a22[6];
					282:word <= a22[7];
					281:word <= a22[8];
					280:word <= a22[9];
					279:word <= a22[10];
					278:word <= a22[11];
					277:word <= a22[12];
					276:word <= a22[13];
					275:word <= a22[14];
					274:word <= a22[15];
					273:word <= a22[16];
					272:word <= a22[17];
					271:word <= a22[18];
					270:word <= a22[19];
					269:word <= a22[20];
					268:word <= a22[21];
					267:word <= a22[22];
					266:word <= a22[23];
					265:word <= a22[24];
					264:word <= a22[25];
					263:word <= a22[26];
					262:word <= a22[27];
					261:word <= a22[28];
					260:word <= a22[29];
					259:word <= a22[30];
					258:word <= a22[31];
					257:word <= a22[32];
					256:word <= a22[33];
					255:word <= a22[34];
					254:word <= a22[35];
					253:word <= a22[36];
					252:word <= a22[37];
					251:word <= a22[38];
					250:word <= a22[39];
					249:word <= a22[40];
					248:word <= a22[41];
					247:word <= a22[42];
					246:word <= a22[43];
					245:word <= a22[44];
					244:word <= a22[45];
					243:word <= a22[46];
					242:word <= a22[47];
					241:word <= a22[48];
					240:word <= a22[49];
					239:word <= a22[50];
					238:word <= a22[51];
					237:word <= a22[52];
					236:word <= a22[53];
					235:word <= a22[54];
					234:word <= a22[55];
					233:word <= a22[56];
					232:word <= a22[57];
					231:word <= a22[58];
					230:word <= a22[59];
					229:word <= a22[60];
					228:word <= a22[61];
					227:word <= a22[62];
					226:word <= a22[63];
					225:word <= a22[64];
					224:word <= a22[65];
					223:word <= a22[66];
					222:word <= a22[67];
					221:word <= a22[68];
					220:word <= a22[69];
					219:word <= a22[70];
					218:word <= a22[71];
					217:word <= a22[72];
					216:word <= a22[73];
					215:word <= a22[74];
					214:word <= a22[75];
					213:word <= a22[76];
					212:word <= a22[77];
					211:word <= a22[78];
					default:word <= a22[79];
					endcase
				end
				63:begin
				case(x)
					290:word <= a23[0];
					289:word <= a23[1];
					287:word <= a23[2];
					286:word <= a23[3];
					285:word <= a23[4];
					284:word <= a23[5];
					283:word <= a23[6];
					282:word <= a23[7];
					281:word <= a23[8];
					280:word <= a23[9];
					279:word <= a23[10];
					278:word <= a23[11];
					277:word <= a23[12];
					276:word <= a23[13];
					275:word <= a23[14];
					274:word <= a23[15];
					273:word <= a23[16];
					272:word <= a23[17];
					271:word <= a23[18];
					270:word <= a23[19];
					269:word <= a23[20];
					268:word <= a23[21];
					267:word <= a23[22];
					266:word <= a23[23];
					265:word <= a23[24];
					264:word <= a23[25];
					263:word <= a23[26];
					262:word <= a23[27];
					261:word <= a23[28];
					260:word <= a23[29];
					259:word <= a23[30];
					258:word <= a23[31];
					257:word <= a23[32];
					256:word <= a23[33];
					255:word <= a23[34];
					254:word <= a23[35];
					253:word <= a23[36];
					252:word <= a23[37];
					251:word <= a23[38];
					250:word <= a23[39];
					249:word <= a23[40];
					248:word <= a23[41];
					247:word <= a23[42];
					246:word <= a23[43];
					245:word <= a23[44];
					244:word <= a23[45];
					243:word <= a23[46];
					242:word <= a23[47];
					241:word <= a23[48];
					240:word <= a23[49];
					239:word <= a23[50];
					238:word <= a23[51];
					237:word <= a23[52];
					236:word <= a23[53];
					235:word <= a23[54];
					234:word <= a23[55];
					233:word <= a23[56];
					232:word <= a23[57];
					231:word <= a23[58];
					230:word <= a23[59];
					229:word <= a23[60];
					228:word <= a23[61];
					227:word <= a23[62];
					226:word <= a23[63];
					225:word <= a23[64];
					224:word <= a23[65];
					223:word <= a23[66];
					222:word <= a23[67];
					221:word <= a23[68];
					220:word <= a23[69];
					219:word <= a23[70];
					218:word <= a23[71];
					217:word <= a23[72];
					216:word <= a23[73];
					215:word <= a23[74];
					214:word <= a23[75];
					213:word <= a23[76];
					212:word <= a23[77];
					211:word <= a23[78];
					default:word <= a23[79];
					endcase
				end
				64:begin
				case(x)
					290:word <= a24[0];
					289:word <= a24[1];
					287:word <= a24[2];
					286:word <= a24[3];
					285:word <= a24[4];
					284:word <= a24[5];
					283:word <= a24[6];
					282:word <= a24[7];
					281:word <= a24[8];
					280:word <= a24[9];
					279:word <= a24[10];
					278:word <= a24[11];
					277:word <= a24[12];
					276:word <= a24[13];
					275:word <= a24[14];
					274:word <= a24[15];
					273:word <= a24[16];
					272:word <= a24[17];
					271:word <= a24[18];
					270:word <= a24[19];
					269:word <= a24[20];
					268:word <= a24[21];
					267:word <= a24[22];
					266:word <= a24[23];
					265:word <= a24[24];
					264:word <= a24[25];
					263:word <= a24[26];
					262:word <= a24[27];
					261:word <= a24[28];
					260:word <= a24[29];
					259:word <= a24[30];
					258:word <= a24[31];
					257:word <= a24[32];
					256:word <= a24[33];
					255:word <= a24[34];
					254:word <= a24[35];
					253:word <= a24[36];
					252:word <= a24[37];
					251:word <= a24[38];
					250:word <= a24[39];
					249:word <= a24[40];
					248:word <= a24[41];
					247:word <= a24[42];
					246:word <= a24[43];
					245:word <= a24[44];
					244:word <= a24[45];
					243:word <= a24[46];
					242:word <= a24[47];
					241:word <= a24[48];
					240:word <= a24[49];
					239:word <= a24[50];
					238:word <= a24[51];
					237:word <= a24[52];
					236:word <= a24[53];
					235:word <= a24[54];
					234:word <= a24[55];
					233:word <= a24[56];
					232:word <= a24[57];
					231:word <= a24[58];
					230:word <= a24[59];
					229:word <= a24[60];
					228:word <= a24[61];
					227:word <= a24[62];
					226:word <= a24[63];
					225:word <= a24[64];
					224:word <= a24[65];
					223:word <= a24[66];
					222:word <= a24[67];
					221:word <= a24[68];
					220:word <= a24[69];
					219:word <= a24[70];
					218:word <= a24[71];
					217:word <= a24[72];
					216:word <= a24[73];
					215:word <= a24[74];
					214:word <= a24[75];
					213:word <= a24[76];
					212:word <= a24[77];
					211:word <= a24[78];
					default:word <= a24[79];
					endcase
				end
				65:begin
				case(x)
					290:word <= a25[0];
					289:word <= a25[1];
					287:word <= a25[2];
					286:word <= a25[3];
					285:word <= a25[4];
					284:word <= a25[5];
					283:word <= a25[6];
					282:word <= a25[7];
					281:word <= a25[8];
					280:word <= a25[9];
					279:word <= a25[10];
					278:word <= a25[11];
					277:word <= a25[12];
					276:word <= a25[13];
					275:word <= a25[14];
					274:word <= a25[15];
					273:word <= a25[16];
					272:word <= a25[17];
					271:word <= a25[18];
					270:word <= a25[19];
					269:word <= a25[20];
					268:word <= a25[21];
					267:word <= a25[22];
					266:word <= a25[23];
					265:word <= a25[24];
					264:word <= a25[25];
					263:word <= a25[26];
					262:word <= a25[27];
					261:word <= a25[28];
					260:word <= a25[29];
					259:word <= a25[30];
					258:word <= a25[31];
					257:word <= a25[32];
					256:word <= a25[33];
					255:word <= a25[34];
					254:word <= a25[35];
					253:word <= a25[36];
					252:word <= a25[37];
					251:word <= a25[38];
					250:word <= a25[39];
					249:word <= a25[40];
					248:word <= a25[41];
					247:word <= a25[42];
					246:word <= a25[43];
					245:word <= a25[44];
					244:word <= a25[45];
					243:word <= a25[46];
					242:word <= a25[47];
					241:word <= a25[48];
					240:word <= a25[49];
					239:word <= a25[50];
					238:word <= a25[51];
					237:word <= a25[52];
					236:word <= a25[53];
					235:word <= a25[54];
					234:word <= a25[55];
					233:word <= a25[56];
					232:word <= a25[57];
					231:word <= a25[58];
					230:word <= a25[59];
					229:word <= a25[60];
					228:word <= a25[61];
					227:word <= a25[62];
					226:word <= a25[63];
					225:word <= a25[64];
					224:word <= a25[65];
					223:word <= a25[66];
					222:word <= a25[67];
					221:word <= a25[68];
					220:word <= a25[69];
					219:word <= a25[70];
					218:word <= a25[71];
					217:word <= a25[72];
					216:word <= a25[73];
					215:word <= a25[74];
					214:word <= a25[75];
					213:word <= a25[76];
					212:word <= a25[77];
					211:word <= a25[78];
					default:word <= a25[79];
					endcase
				end
				66:begin
				case(x)
					290:word <= a26[0];
					289:word <= a26[1];
					287:word <= a26[2];
					286:word <= a26[3];
					285:word <= a26[4];
					284:word <= a26[5];
					283:word <= a26[6];
					282:word <= a26[7];
					281:word <= a26[8];
					280:word <= a26[9];
					279:word <= a26[10];
					278:word <= a26[11];
					277:word <= a26[12];
					276:word <= a26[13];
					275:word <= a26[14];
					274:word <= a26[15];
					273:word <= a26[16];
					272:word <= a26[17];
					271:word <= a26[18];
					270:word <= a26[19];
					269:word <= a26[20];
					268:word <= a26[21];
					267:word <= a26[22];
					266:word <= a26[23];
					265:word <= a26[24];
					264:word <= a26[25];
					263:word <= a26[26];
					262:word <= a26[27];
					261:word <= a26[28];
					260:word <= a26[29];
					259:word <= a26[30];
					258:word <= a26[31];
					257:word <= a26[32];
					256:word <= a26[33];
					255:word <= a26[34];
					254:word <= a26[35];
					253:word <= a26[36];
					252:word <= a26[37];
					251:word <= a26[38];
					250:word <= a26[39];
					249:word <= a26[40];
					248:word <= a26[41];
					247:word <= a26[42];
					246:word <= a26[43];
					245:word <= a26[44];
					244:word <= a26[45];
					243:word <= a26[46];
					242:word <= a26[47];
					241:word <= a26[48];
					240:word <= a26[49];
					239:word <= a26[50];
					238:word <= a26[51];
					237:word <= a26[52];
					236:word <= a26[53];
					235:word <= a26[54];
					234:word <= a26[55];
					233:word <= a26[56];
					232:word <= a26[57];
					231:word <= a26[58];
					230:word <= a26[59];
					229:word <= a26[60];
					228:word <= a26[61];
					227:word <= a26[62];
					226:word <= a26[63];
					225:word <= a26[64];
					224:word <= a26[65];
					223:word <= a26[66];
					222:word <= a26[67];
					221:word <= a26[68];
					220:word <= a26[69];
					219:word <= a26[70];
					218:word <= a26[71];
					217:word <= a26[72];
					216:word <= a26[73];
					215:word <= a26[74];
					214:word <= a26[75];
					213:word <= a26[76];
					212:word <= a26[77];
					211:word <= a26[78];
					default:word <= a26[79];
					endcase
				end
				67:begin
				case(x)
					290:word <= a27[0];
					289:word <= a27[1];
					287:word <= a27[2];
					286:word <= a27[3];
					285:word <= a27[4];
					284:word <= a27[5];
					283:word <= a27[6];
					282:word <= a27[7];
					281:word <= a27[8];
					280:word <= a27[9];
					279:word <= a27[10];
					278:word <= a27[11];
					277:word <= a27[12];
					276:word <= a27[13];
					275:word <= a27[14];
					274:word <= a27[15];
					273:word <= a27[16];
					272:word <= a27[17];
					271:word <= a27[18];
					270:word <= a27[19];
					269:word <= a27[20];
					268:word <= a27[21];
					267:word <= a27[22];
					266:word <= a27[23];
					265:word <= a27[24];
					264:word <= a27[25];
					263:word <= a27[26];
					262:word <= a27[27];
					261:word <= a27[28];
					260:word <= a27[29];
					259:word <= a27[30];
					258:word <= a27[31];
					257:word <= a27[32];
					256:word <= a27[33];
					255:word <= a27[34];
					254:word <= a27[35];
					253:word <= a27[36];
					252:word <= a27[37];
					251:word <= a27[38];
					250:word <= a27[39];
					249:word <= a27[40];
					248:word <= a27[41];
					247:word <= a27[42];
					246:word <= a27[43];
					245:word <= a27[44];
					244:word <= a27[45];
					243:word <= a27[46];
					242:word <= a27[47];
					241:word <= a27[48];
					240:word <= a27[49];
					239:word <= a27[50];
					238:word <= a27[51];
					237:word <= a27[52];
					236:word <= a27[53];
					235:word <= a27[54];
					234:word <= a27[55];
					233:word <= a27[56];
					232:word <= a27[57];
					231:word <= a27[58];
					230:word <= a27[59];
					229:word <= a27[60];
					228:word <= a27[61];
					227:word <= a27[62];
					226:word <= a27[63];
					225:word <= a27[64];
					224:word <= a27[65];
					223:word <= a27[66];
					222:word <= a27[67];
					221:word <= a27[68];
					220:word <= a27[69];
					219:word <= a27[70];
					218:word <= a27[71];
					217:word <= a27[72];
					216:word <= a27[73];
					215:word <= a27[74];
					214:word <= a27[75];
					213:word <= a27[76];
					212:word <= a27[77];
					211:word <= a27[78];
					default:word <= a27[79];
					endcase
				end
				68:begin
				case(x)
					290:word <= a28[0];
					289:word <= a28[1];
					287:word <= a28[2];
					286:word <= a28[3];
					285:word <= a28[4];
					284:word <= a28[5];
					283:word <= a28[6];
					282:word <= a28[7];
					281:word <= a28[8];
					280:word <= a28[9];
					279:word <= a28[10];
					278:word <= a28[11];
					277:word <= a28[12];
					276:word <= a28[13];
					275:word <= a28[14];
					274:word <= a28[15];
					273:word <= a28[16];
					272:word <= a28[17];
					271:word <= a28[18];
					270:word <= a28[19];
					269:word <= a28[20];
					268:word <= a28[21];
					267:word <= a28[22];
					266:word <= a28[23];
					265:word <= a28[24];
					264:word <= a28[25];
					263:word <= a28[26];
					262:word <= a28[27];
					261:word <= a28[28];
					260:word <= a28[29];
					259:word <= a28[30];
					258:word <= a28[31];
					257:word <= a28[32];
					256:word <= a28[33];
					255:word <= a28[34];
					254:word <= a28[35];
					253:word <= a28[36];
					252:word <= a28[37];
					251:word <= a28[38];
					250:word <= a28[39];
					249:word <= a28[40];
					248:word <= a28[41];
					247:word <= a28[42];
					246:word <= a28[43];
					245:word <= a28[44];
					244:word <= a28[45];
					243:word <= a28[46];
					242:word <= a28[47];
					241:word <= a28[48];
					240:word <= a28[49];
					239:word <= a28[50];
					238:word <= a28[51];
					237:word <= a28[52];
					236:word <= a28[53];
					235:word <= a28[54];
					234:word <= a28[55];
					233:word <= a28[56];
					232:word <= a28[57];
					231:word <= a28[58];
					230:word <= a28[59];
					229:word <= a28[60];
					228:word <= a28[61];
					227:word <= a28[62];
					226:word <= a28[63];
					225:word <= a28[64];
					224:word <= a28[65];
					223:word <= a28[66];
					222:word <= a28[67];
					221:word <= a28[68];
					220:word <= a28[69];
					219:word <= a28[70];
					218:word <= a28[71];
					217:word <= a28[72];
					216:word <= a28[73];
					215:word <= a28[74];
					214:word <= a28[75];
					213:word <= a28[76];
					212:word <= a28[77];
					211:word <= a28[78];
					default:word <= a28[79];
					endcase
				end
				69:begin
				case(x)
					290:word <= a29[0];
					289:word <= a29[1];
					287:word <= a29[2];
					286:word <= a29[3];
					285:word <= a29[4];
					284:word <= a29[5];
					283:word <= a29[6];
					282:word <= a29[7];
					281:word <= a29[8];
					280:word <= a29[9];
					279:word <= a29[10];
					278:word <= a29[11];
					277:word <= a29[12];
					276:word <= a29[13];
					275:word <= a29[14];
					274:word <= a29[15];
					273:word <= a29[16];
					272:word <= a29[17];
					271:word <= a29[18];
					270:word <= a29[19];
					269:word <= a29[20];
					268:word <= a29[21];
					267:word <= a29[22];
					266:word <= a29[23];
					265:word <= a29[24];
					264:word <= a29[25];
					263:word <= a29[26];
					262:word <= a29[27];
					261:word <= a29[28];
					260:word <= a29[29];
					259:word <= a29[30];
					258:word <= a29[31];
					257:word <= a29[32];
					256:word <= a29[33];
					255:word <= a29[34];
					254:word <= a29[35];
					253:word <= a29[36];
					252:word <= a29[37];
					251:word <= a29[38];
					250:word <= a29[39];
					249:word <= a29[40];
					248:word <= a29[41];
					247:word <= a29[42];
					246:word <= a29[43];
					245:word <= a29[44];
					244:word <= a29[45];
					243:word <= a29[46];
					242:word <= a29[47];
					241:word <= a29[48];
					240:word <= a29[49];
					239:word <= a29[50];
					238:word <= a29[51];
					237:word <= a29[52];
					236:word <= a29[53];
					235:word <= a29[54];
					234:word <= a29[55];
					233:word <= a29[56];
					232:word <= a29[57];
					231:word <= a29[58];
					230:word <= a29[59];
					229:word <= a29[60];
					228:word <= a29[61];
					227:word <= a29[62];
					226:word <= a29[63];
					225:word <= a29[64];
					224:word <= a29[65];
					223:word <= a29[66];
					222:word <= a29[67];
					221:word <= a29[68];
					220:word <= a29[69];
					219:word <= a29[70];
					218:word <= a29[71];
					217:word <= a29[72];
					216:word <= a29[73];
					215:word <= a29[74];
					214:word <= a29[75];
					213:word <= a29[76];
					212:word <= a29[77];
					211:word <= a29[78];
					default:word <= a29[79];
					endcase
				end
				70:begin
				case(x)
					290:word <= a30[0];
					289:word <= a30[1];
					287:word <= a30[2];
					286:word <= a30[3];
					285:word <= a30[4];
					284:word <= a30[5];
					283:word <= a30[6];
					282:word <= a30[7];
					281:word <= a30[8];
					280:word <= a30[9];
					279:word <= a30[10];
					278:word <= a30[11];
					277:word <= a30[12];
					276:word <= a30[13];
					275:word <= a30[14];
					274:word <= a30[15];
					273:word <= a30[16];
					272:word <= a30[17];
					271:word <= a30[18];
					270:word <= a30[19];
					269:word <= a30[20];
					268:word <= a30[21];
					267:word <= a30[22];
					266:word <= a30[23];
					265:word <= a30[24];
					264:word <= a30[25];
					263:word <= a30[26];
					262:word <= a30[27];
					261:word <= a30[28];
					260:word <= a30[29];
					259:word <= a30[30];
					258:word <= a30[31];
					257:word <= a30[32];
					256:word <= a30[33];
					255:word <= a30[34];
					254:word <= a30[35];
					253:word <= a30[36];
					252:word <= a30[37];
					251:word <= a30[38];
					250:word <= a30[39];
					249:word <= a30[40];
					248:word <= a30[41];
					247:word <= a30[42];
					246:word <= a30[43];
					245:word <= a30[44];
					244:word <= a30[45];
					243:word <= a30[46];
					242:word <= a30[47];
					241:word <= a30[48];
					240:word <= a30[49];
					239:word <= a30[50];
					238:word <= a30[51];
					237:word <= a30[52];
					236:word <= a30[53];
					235:word <= a30[54];
					234:word <= a30[55];
					233:word <= a30[56];
					232:word <= a30[57];
					231:word <= a30[58];
					230:word <= a30[59];
					229:word <= a30[60];
					228:word <= a30[61];
					227:word <= a30[62];
					226:word <= a30[63];
					225:word <= a30[64];
					224:word <= a30[65];
					223:word <= a30[66];
					222:word <= a30[67];
					221:word <= a30[68];
					220:word <= a30[69];
					219:word <= a30[70];
					218:word <= a30[71];
					217:word <= a30[72];
					216:word <= a30[73];
					215:word <= a30[74];
					214:word <= a30[75];
					213:word <= a30[76];
					212:word <= a30[77];
					211:word <= a30[78];
					default:word <= a30[79];
					endcase
				end
				71:begin
				case(x)
					290:word <= a31[0];
					289:word <= a31[1];
					287:word <= a31[2];
					286:word <= a31[3];
					285:word <= a31[4];
					284:word <= a31[5];
					283:word <= a31[6];
					282:word <= a31[7];
					281:word <= a31[8];
					280:word <= a31[9];
					279:word <= a31[10];
					278:word <= a31[11];
					277:word <= a31[12];
					276:word <= a31[13];
					275:word <= a31[14];
					274:word <= a31[15];
					273:word <= a31[16];
					272:word <= a31[17];
					271:word <= a31[18];
					270:word <= a31[19];
					269:word <= a31[20];
					268:word <= a31[21];
					267:word <= a31[22];
					266:word <= a31[23];
					265:word <= a31[24];
					264:word <= a31[25];
					263:word <= a31[26];
					262:word <= a31[27];
					261:word <= a31[28];
					260:word <= a31[29];
					259:word <= a31[30];
					258:word <= a31[31];
					257:word <= a31[32];
					256:word <= a31[33];
					255:word <= a31[34];
					254:word <= a31[35];
					253:word <= a31[36];
					252:word <= a31[37];
					251:word <= a31[38];
					250:word <= a31[39];
					249:word <= a31[40];
					248:word <= a31[41];
					247:word <= a31[42];
					246:word <= a31[43];
					245:word <= a31[44];
					244:word <= a31[45];
					243:word <= a31[46];
					242:word <= a31[47];
					241:word <= a31[48];
					240:word <= a31[49];
					239:word <= a31[50];
					238:word <= a31[51];
					237:word <= a31[52];
					236:word <= a31[53];
					235:word <= a31[54];
					234:word <= a31[55];
					233:word <= a31[56];
					232:word <= a31[57];
					231:word <= a31[58];
					230:word <= a31[59];
					229:word <= a31[60];
					228:word <= a31[61];
					227:word <= a31[62];
					226:word <= a31[63];
					225:word <= a31[64];
					224:word <= a31[65];
					223:word <= a31[66];
					222:word <= a31[67];
					221:word <= a31[68];
					220:word <= a31[69];
					219:word <= a31[70];
					218:word <= a31[71];
					217:word <= a31[72];
					216:word <= a31[73];
					215:word <= a31[74];
					214:word <= a31[75];
					213:word <= a31[76];
					212:word <= a31[77];
					211:word <= a31[78];
					default:word <= a31[79];
					endcase
				end
				72:begin
				case(x)
					290:word <= a32[0];
					289:word <= a32[1];
					287:word <= a32[2];
					286:word <= a32[3];
					285:word <= a32[4];
					284:word <= a32[5];
					283:word <= a32[6];
					282:word <= a32[7];
					281:word <= a32[8];
					280:word <= a32[9];
					279:word <= a32[10];
					278:word <= a32[11];
					277:word <= a32[12];
					276:word <= a32[13];
					275:word <= a32[14];
					274:word <= a32[15];
					273:word <= a32[16];
					272:word <= a32[17];
					271:word <= a32[18];
					270:word <= a32[19];
					269:word <= a32[20];
					268:word <= a32[21];
					267:word <= a32[22];
					266:word <= a32[23];
					265:word <= a32[24];
					264:word <= a32[25];
					263:word <= a32[26];
					262:word <= a32[27];
					261:word <= a32[28];
					260:word <= a32[29];
					259:word <= a32[30];
					258:word <= a32[31];
					257:word <= a32[32];
					256:word <= a32[33];
					255:word <= a32[34];
					254:word <= a32[35];
					253:word <= a32[36];
					252:word <= a32[37];
					251:word <= a32[38];
					250:word <= a32[39];
					249:word <= a32[40];
					248:word <= a32[41];
					247:word <= a32[42];
					246:word <= a32[43];
					245:word <= a32[44];
					244:word <= a32[45];
					243:word <= a32[46];
					242:word <= a32[47];
					241:word <= a32[48];
					240:word <= a32[49];
					239:word <= a32[50];
					238:word <= a32[51];
					237:word <= a32[52];
					236:word <= a32[53];
					235:word <= a32[54];
					234:word <= a32[55];
					233:word <= a32[56];
					232:word <= a32[57];
					231:word <= a32[58];
					230:word <= a32[59];
					229:word <= a32[60];
					228:word <= a32[61];
					227:word <= a32[62];
					226:word <= a32[63];
					225:word <= a32[64];
					224:word <= a32[65];
					223:word <= a32[66];
					222:word <= a32[67];
					221:word <= a32[68];
					220:word <= a32[69];
					219:word <= a32[70];
					218:word <= a32[71];
					217:word <= a32[72];
					216:word <= a32[73];
					215:word <= a32[74];
					214:word <= a32[75];
					213:word <= a32[76];
					212:word <= a32[77];
					211:word <= a32[78];
					default:word <= a32[79];
					endcase
				end
				73:begin
				case(x)
					290:word <= a33[0];
					289:word <= a33[1];
					287:word <= a33[2];
					286:word <= a33[3];
					285:word <= a33[4];
					284:word <= a33[5];
					283:word <= a33[6];
					282:word <= a33[7];
					281:word <= a33[8];
					280:word <= a33[9];
					279:word <= a33[10];
					278:word <= a33[11];
					277:word <= a33[12];
					276:word <= a33[13];
					275:word <= a33[14];
					274:word <= a33[15];
					273:word <= a33[16];
					272:word <= a33[17];
					271:word <= a33[18];
					270:word <= a33[19];
					269:word <= a33[20];
					268:word <= a33[21];
					267:word <= a33[22];
					266:word <= a33[23];
					265:word <= a33[24];
					264:word <= a33[25];
					263:word <= a33[26];
					262:word <= a33[27];
					261:word <= a33[28];
					260:word <= a33[29];
					259:word <= a33[30];
					258:word <= a33[31];
					257:word <= a33[32];
					256:word <= a33[33];
					255:word <= a33[34];
					254:word <= a33[35];
					253:word <= a33[36];
					252:word <= a33[37];
					251:word <= a33[38];
					250:word <= a33[39];
					249:word <= a33[40];
					248:word <= a33[41];
					247:word <= a33[42];
					246:word <= a33[43];
					245:word <= a33[44];
					244:word <= a33[45];
					243:word <= a33[46];
					242:word <= a33[47];
					241:word <= a33[48];
					240:word <= a33[49];
					239:word <= a33[50];
					238:word <= a33[51];
					237:word <= a33[52];
					236:word <= a33[53];
					235:word <= a33[54];
					234:word <= a33[55];
					233:word <= a33[56];
					232:word <= a33[57];
					231:word <= a33[58];
					230:word <= a33[59];
					229:word <= a33[60];
					228:word <= a33[61];
					227:word <= a33[62];
					226:word <= a33[63];
					225:word <= a33[64];
					224:word <= a33[65];
					223:word <= a33[66];
					222:word <= a33[67];
					221:word <= a33[68];
					220:word <= a33[69];
					219:word <= a33[70];
					218:word <= a33[71];
					217:word <= a33[72];
					216:word <= a33[73];
					215:word <= a33[74];
					214:word <= a33[75];
					213:word <= a33[76];
					212:word <= a33[77];
					211:word <= a33[78];
					default:word <= a33[79];
					endcase
				end
				74:begin
				case(x)
					290:word <= a34[0];
					289:word <= a34[1];
					287:word <= a34[2];
					286:word <= a34[3];
					285:word <= a34[4];
					284:word <= a34[5];
					283:word <= a34[6];
					282:word <= a34[7];
					281:word <= a34[8];
					280:word <= a34[9];
					279:word <= a34[10];
					278:word <= a34[11];
					277:word <= a34[12];
					276:word <= a34[13];
					275:word <= a34[14];
					274:word <= a34[15];
					273:word <= a34[16];
					272:word <= a34[17];
					271:word <= a34[18];
					270:word <= a34[19];
					269:word <= a34[20];
					268:word <= a34[21];
					267:word <= a34[22];
					266:word <= a34[23];
					265:word <= a34[24];
					264:word <= a34[25];
					263:word <= a34[26];
					262:word <= a34[27];
					261:word <= a34[28];
					260:word <= a34[29];
					259:word <= a34[30];
					258:word <= a34[31];
					257:word <= a34[32];
					256:word <= a34[33];
					255:word <= a34[34];
					254:word <= a34[35];
					253:word <= a34[36];
					252:word <= a34[37];
					251:word <= a34[38];
					250:word <= a34[39];
					249:word <= a34[40];
					248:word <= a34[41];
					247:word <= a34[42];
					246:word <= a34[43];
					245:word <= a34[44];
					244:word <= a34[45];
					243:word <= a34[46];
					242:word <= a34[47];
					241:word <= a34[48];
					240:word <= a34[49];
					239:word <= a34[50];
					238:word <= a34[51];
					237:word <= a34[52];
					236:word <= a34[53];
					235:word <= a34[54];
					234:word <= a34[55];
					233:word <= a34[56];
					232:word <= a34[57];
					231:word <= a34[58];
					230:word <= a34[59];
					229:word <= a34[60];
					228:word <= a34[61];
					227:word <= a34[62];
					226:word <= a34[63];
					225:word <= a34[64];
					224:word <= a34[65];
					223:word <= a34[66];
					222:word <= a34[67];
					221:word <= a34[68];
					220:word <= a34[69];
					219:word <= a34[70];
					218:word <= a34[71];
					217:word <= a34[72];
					216:word <= a34[73];
					215:word <= a34[74];
					214:word <= a34[75];
					213:word <= a34[76];
					212:word <= a34[77];
					211:word <= a34[78];
					default:word <= a34[79];
					endcase
				end
				75:begin
				case(x)
					290:word <= a35[0];
					289:word <= a35[1];
					287:word <= a35[2];
					286:word <= a35[3];
					285:word <= a35[4];
					284:word <= a35[5];
					283:word <= a35[6];
					282:word <= a35[7];
					281:word <= a35[8];
					280:word <= a35[9];
					279:word <= a35[10];
					278:word <= a35[11];
					277:word <= a35[12];
					276:word <= a35[13];
					275:word <= a35[14];
					274:word <= a35[15];
					273:word <= a35[16];
					272:word <= a35[17];
					271:word <= a35[18];
					270:word <= a35[19];
					269:word <= a35[20];
					268:word <= a35[21];
					267:word <= a35[22];
					266:word <= a35[23];
					265:word <= a35[24];
					264:word <= a35[25];
					263:word <= a35[26];
					262:word <= a35[27];
					261:word <= a35[28];
					260:word <= a35[29];
					259:word <= a35[30];
					258:word <= a35[31];
					257:word <= a35[32];
					256:word <= a35[33];
					255:word <= a35[34];
					254:word <= a35[35];
					253:word <= a35[36];
					252:word <= a35[37];
					251:word <= a35[38];
					250:word <= a35[39];
					249:word <= a35[40];
					248:word <= a35[41];
					247:word <= a35[42];
					246:word <= a35[43];
					245:word <= a35[44];
					244:word <= a35[45];
					243:word <= a35[46];
					242:word <= a35[47];
					241:word <= a35[48];
					240:word <= a35[49];
					239:word <= a35[50];
					238:word <= a35[51];
					237:word <= a35[52];
					236:word <= a35[53];
					235:word <= a35[54];
					234:word <= a35[55];
					233:word <= a35[56];
					232:word <= a35[57];
					231:word <= a35[58];
					230:word <= a35[59];
					229:word <= a35[60];
					228:word <= a35[61];
					227:word <= a35[62];
					226:word <= a35[63];
					225:word <= a35[64];
					224:word <= a35[65];
					223:word <= a35[66];
					222:word <= a35[67];
					221:word <= a35[68];
					220:word <= a35[69];
					219:word <= a35[70];
					218:word <= a35[71];
					217:word <= a35[72];
					216:word <= a35[73];
					215:word <= a35[74];
					214:word <= a35[75];
					213:word <= a35[76];
					212:word <= a35[77];
					211:word <= a35[78];
					default:word <= a35[79];
					endcase
				end
				76:begin
				case(x)
					290:word <= a36[0];
					289:word <= a36[1];
					287:word <= a36[2];
					286:word <= a36[3];
					285:word <= a36[4];
					284:word <= a36[5];
					283:word <= a36[6];
					282:word <= a36[7];
					281:word <= a36[8];
					280:word <= a36[9];
					279:word <= a36[10];
					278:word <= a36[11];
					277:word <= a36[12];
					276:word <= a36[13];
					275:word <= a36[14];
					274:word <= a36[15];
					273:word <= a36[16];
					272:word <= a36[17];
					271:word <= a36[18];
					270:word <= a36[19];
					269:word <= a36[20];
					268:word <= a36[21];
					267:word <= a36[22];
					266:word <= a36[23];
					265:word <= a36[24];
					264:word <= a36[25];
					263:word <= a36[26];
					262:word <= a36[27];
					261:word <= a36[28];
					260:word <= a36[29];
					259:word <= a36[30];
					258:word <= a36[31];
					257:word <= a36[32];
					256:word <= a36[33];
					255:word <= a36[34];
					254:word <= a36[35];
					253:word <= a36[36];
					252:word <= a36[37];
					251:word <= a36[38];
					250:word <= a36[39];
					249:word <= a36[40];
					248:word <= a36[41];
					247:word <= a36[42];
					246:word <= a36[43];
					245:word <= a36[44];
					244:word <= a36[45];
					243:word <= a36[46];
					242:word <= a36[47];
					241:word <= a36[48];
					240:word <= a36[49];
					239:word <= a36[50];
					238:word <= a36[51];
					237:word <= a36[52];
					236:word <= a36[53];
					235:word <= a36[54];
					234:word <= a36[55];
					233:word <= a36[56];
					232:word <= a36[57];
					231:word <= a36[58];
					230:word <= a36[59];
					229:word <= a36[60];
					228:word <= a36[61];
					227:word <= a36[62];
					226:word <= a36[63];
					225:word <= a36[64];
					224:word <= a36[65];
					223:word <= a36[66];
					222:word <= a36[67];
					221:word <= a36[68];
					220:word <= a36[69];
					219:word <= a36[70];
					218:word <= a36[71];
					217:word <= a36[72];
					216:word <= a36[73];
					215:word <= a36[74];
					214:word <= a36[75];
					213:word <= a36[76];
					212:word <= a36[77];
					211:word <= a36[78];
					default:word <= a36[79];
					endcase
				end
				77:begin
				case(x)
					290:word <= a37[0];
					289:word <= a37[1];
					287:word <= a37[2];
					286:word <= a37[3];
					285:word <= a37[4];
					284:word <= a37[5];
					283:word <= a37[6];
					282:word <= a37[7];
					281:word <= a37[8];
					280:word <= a37[9];
					279:word <= a37[10];
					278:word <= a37[11];
					277:word <= a37[12];
					276:word <= a37[13];
					275:word <= a37[14];
					274:word <= a37[15];
					273:word <= a37[16];
					272:word <= a37[17];
					271:word <= a37[18];
					270:word <= a37[19];
					269:word <= a37[20];
					268:word <= a37[21];
					267:word <= a37[22];
					266:word <= a37[23];
					265:word <= a37[24];
					264:word <= a37[25];
					263:word <= a37[26];
					262:word <= a37[27];
					261:word <= a37[28];
					260:word <= a37[29];
					259:word <= a37[30];
					258:word <= a37[31];
					257:word <= a37[32];
					256:word <= a37[33];
					255:word <= a37[34];
					254:word <= a37[35];
					253:word <= a37[36];
					252:word <= a37[37];
					251:word <= a37[38];
					250:word <= a37[39];
					249:word <= a37[40];
					248:word <= a37[41];
					247:word <= a37[42];
					246:word <= a37[43];
					245:word <= a37[44];
					244:word <= a37[45];
					243:word <= a37[46];
					242:word <= a37[47];
					241:word <= a37[48];
					240:word <= a37[49];
					239:word <= a37[50];
					238:word <= a37[51];
					237:word <= a37[52];
					236:word <= a37[53];
					235:word <= a37[54];
					234:word <= a37[55];
					233:word <= a37[56];
					232:word <= a37[57];
					231:word <= a37[58];
					230:word <= a37[59];
					229:word <= a37[60];
					228:word <= a37[61];
					227:word <= a37[62];
					226:word <= a37[63];
					225:word <= a37[64];
					224:word <= a37[65];
					223:word <= a37[66];
					222:word <= a37[67];
					221:word <= a37[68];
					220:word <= a37[69];
					219:word <= a37[70];
					218:word <= a37[71];
					217:word <= a37[72];
					216:word <= a37[73];
					215:word <= a37[74];
					214:word <= a37[75];
					213:word <= a37[76];
					212:word <= a37[77];
					211:word <= a37[78];
					default:word <= a37[79];
					endcase
				end
				78:begin
				case(x)
					290:word <= a38[0];
					289:word <= a38[1];
					287:word <= a38[2];
					286:word <= a38[3];
					285:word <= a38[4];
					284:word <= a38[5];
					283:word <= a38[6];
					282:word <= a38[7];
					281:word <= a38[8];
					280:word <= a38[9];
					279:word <= a38[10];
					278:word <= a38[11];
					277:word <= a38[12];
					276:word <= a38[13];
					275:word <= a38[14];
					274:word <= a38[15];
					273:word <= a38[16];
					272:word <= a38[17];
					271:word <= a38[18];
					270:word <= a38[19];
					269:word <= a38[20];
					268:word <= a38[21];
					267:word <= a38[22];
					266:word <= a38[23];
					265:word <= a38[24];
					264:word <= a38[25];
					263:word <= a38[26];
					262:word <= a38[27];
					261:word <= a38[28];
					260:word <= a38[29];
					259:word <= a38[30];
					258:word <= a38[31];
					257:word <= a38[32];
					256:word <= a38[33];
					255:word <= a38[34];
					254:word <= a38[35];
					253:word <= a38[36];
					252:word <= a38[37];
					251:word <= a38[38];
					250:word <= a38[39];
					249:word <= a38[40];
					248:word <= a38[41];
					247:word <= a38[42];
					246:word <= a38[43];
					245:word <= a38[44];
					244:word <= a38[45];
					243:word <= a38[46];
					242:word <= a38[47];
					241:word <= a38[48];
					240:word <= a38[49];
					239:word <= a38[50];
					238:word <= a38[51];
					237:word <= a38[52];
					236:word <= a38[53];
					235:word <= a38[54];
					234:word <= a38[55];
					233:word <= a38[56];
					232:word <= a38[57];
					231:word <= a38[58];
					230:word <= a38[59];
					229:word <= a38[60];
					228:word <= a38[61];
					227:word <= a38[62];
					226:word <= a38[63];
					225:word <= a38[64];
					224:word <= a38[65];
					223:word <= a38[66];
					222:word <= a38[67];
					221:word <= a38[68];
					220:word <= a38[69];
					219:word <= a38[70];
					218:word <= a38[71];
					217:word <= a38[72];
					216:word <= a38[73];
					215:word <= a38[74];
					214:word <= a38[75];
					213:word <= a38[76];
					212:word <= a38[77];
					211:word <= a38[78];
					default:word <= a38[79];
					endcase
				end
				79:begin
				case(x)
					290:word <= a39[0];
					289:word <= a39[1];
					287:word <= a39[2];
					286:word <= a39[3];
					285:word <= a39[4];
					284:word <= a39[5];
					283:word <= a39[6];
					282:word <= a39[7];
					281:word <= a39[8];
					280:word <= a39[9];
					279:word <= a39[10];
					278:word <= a39[11];
					277:word <= a39[12];
					276:word <= a39[13];
					275:word <= a39[14];
					274:word <= a39[15];
					273:word <= a39[16];
					272:word <= a39[17];
					271:word <= a39[18];
					270:word <= a39[19];
					269:word <= a39[20];
					268:word <= a39[21];
					267:word <= a39[22];
					266:word <= a39[23];
					265:word <= a39[24];
					264:word <= a39[25];
					263:word <= a39[26];
					262:word <= a39[27];
					261:word <= a39[28];
					260:word <= a39[29];
					259:word <= a39[30];
					258:word <= a39[31];
					257:word <= a39[32];
					256:word <= a39[33];
					255:word <= a39[34];
					254:word <= a39[35];
					253:word <= a39[36];
					252:word <= a39[37];
					251:word <= a39[38];
					250:word <= a39[39];
					249:word <= a39[40];
					248:word <= a39[41];
					247:word <= a39[42];
					246:word <= a39[43];
					245:word <= a39[44];
					244:word <= a39[45];
					243:word <= a39[46];
					242:word <= a39[47];
					241:word <= a39[48];
					240:word <= a39[49];
					239:word <= a39[50];
					238:word <= a39[51];
					237:word <= a39[52];
					236:word <= a39[53];
					235:word <= a39[54];
					234:word <= a39[55];
					233:word <= a39[56];
					232:word <= a39[57];
					231:word <= a39[58];
					230:word <= a39[59];
					229:word <= a39[60];
					228:word <= a39[61];
					227:word <= a39[62];
					226:word <= a39[63];
					225:word <= a39[64];
					224:word <= a39[65];
					223:word <= a39[66];
					222:word <= a39[67];
					221:word <= a39[68];
					220:word <= a39[69];
					219:word <= a39[70];
					218:word <= a39[71];
					217:word <= a39[72];
					216:word <= a39[73];
					215:word <= a39[74];
					214:word <= a39[75];
					213:word <= a39[76];
					212:word <= a39[77];
					211:word <= a39[78];
					default:word <= a39[79];
					endcase
				end
				80:begin
				case(x)
					290:word <= a40[0];
					289:word <= a40[1];
					287:word <= a40[2];
					286:word <= a40[3];
					285:word <= a40[4];
					284:word <= a40[5];
					283:word <= a40[6];
					282:word <= a40[7];
					281:word <= a40[8];
					280:word <= a40[9];
					279:word <= a40[10];
					278:word <= a40[11];
					277:word <= a40[12];
					276:word <= a40[13];
					275:word <= a40[14];
					274:word <= a40[15];
					273:word <= a40[16];
					272:word <= a40[17];
					271:word <= a40[18];
					270:word <= a40[19];
					269:word <= a40[20];
					268:word <= a40[21];
					267:word <= a40[22];
					266:word <= a40[23];
					265:word <= a40[24];
					264:word <= a40[25];
					263:word <= a40[26];
					262:word <= a40[27];
					261:word <= a40[28];
					260:word <= a40[29];
					259:word <= a40[30];
					258:word <= a40[31];
					257:word <= a40[32];
					256:word <= a40[33];
					255:word <= a40[34];
					254:word <= a40[35];
					253:word <= a40[36];
					252:word <= a40[37];
					251:word <= a40[38];
					250:word <= a40[39];
					249:word <= a40[40];
					248:word <= a40[41];
					247:word <= a40[42];
					246:word <= a40[43];
					245:word <= a40[44];
					244:word <= a40[45];
					243:word <= a40[46];
					242:word <= a40[47];
					241:word <= a40[48];
					240:word <= a40[49];
					239:word <= a40[50];
					238:word <= a40[51];
					237:word <= a40[52];
					236:word <= a40[53];
					235:word <= a40[54];
					234:word <= a40[55];
					233:word <= a40[56];
					232:word <= a40[57];
					231:word <= a40[58];
					230:word <= a40[59];
					229:word <= a40[60];
					228:word <= a40[61];
					227:word <= a40[62];
					226:word <= a40[63];
					225:word <= a40[64];
					224:word <= a40[65];
					223:word <= a40[66];
					222:word <= a40[67];
					221:word <= a40[68];
					220:word <= a40[69];
					219:word <= a40[70];
					218:word <= a40[71];
					217:word <= a40[72];
					216:word <= a40[73];
					215:word <= a40[74];
					214:word <= a40[75];
					213:word <= a40[76];
					212:word <= a40[77];
					211:word <= a40[78];
					default:word <= a40[79];
					endcase
				end
				81:begin
				case(x)
					290:word <= a41[0];
					289:word <= a41[1];
					287:word <= a41[2];
					286:word <= a41[3];
					285:word <= a41[4];
					284:word <= a41[5];
					283:word <= a41[6];
					282:word <= a41[7];
					281:word <= a41[8];
					280:word <= a41[9];
					279:word <= a41[10];
					278:word <= a41[11];
					277:word <= a41[12];
					276:word <= a41[13];
					275:word <= a41[14];
					274:word <= a41[15];
					273:word <= a41[16];
					272:word <= a41[17];
					271:word <= a41[18];
					270:word <= a41[19];
					269:word <= a41[20];
					268:word <= a41[21];
					267:word <= a41[22];
					266:word <= a41[23];
					265:word <= a41[24];
					264:word <= a41[25];
					263:word <= a41[26];
					262:word <= a41[27];
					261:word <= a41[28];
					260:word <= a41[29];
					259:word <= a41[30];
					258:word <= a41[31];
					257:word <= a41[32];
					256:word <= a41[33];
					255:word <= a41[34];
					254:word <= a41[35];
					253:word <= a41[36];
					252:word <= a41[37];
					251:word <= a41[38];
					250:word <= a41[39];
					249:word <= a41[40];
					248:word <= a41[41];
					247:word <= a41[42];
					246:word <= a41[43];
					245:word <= a41[44];
					244:word <= a41[45];
					243:word <= a41[46];
					242:word <= a41[47];
					241:word <= a41[48];
					240:word <= a41[49];
					239:word <= a41[50];
					238:word <= a41[51];
					237:word <= a41[52];
					236:word <= a41[53];
					235:word <= a41[54];
					234:word <= a41[55];
					233:word <= a41[56];
					232:word <= a41[57];
					231:word <= a41[58];
					230:word <= a41[59];
					229:word <= a41[60];
					228:word <= a41[61];
					227:word <= a41[62];
					226:word <= a41[63];
					225:word <= a41[64];
					224:word <= a41[65];
					223:word <= a41[66];
					222:word <= a41[67];
					221:word <= a41[68];
					220:word <= a41[69];
					219:word <= a41[70];
					218:word <= a41[71];
					217:word <= a41[72];
					216:word <= a41[73];
					215:word <= a41[74];
					214:word <= a41[75];
					213:word <= a41[76];
					212:word <= a41[77];
					211:word <= a41[78];
					default:word <= a41[79];
					endcase
				end
				82:begin
				case(x)
					290:word <= a42[0];
					289:word <= a42[1];
					287:word <= a42[2];
					286:word <= a42[3];
					285:word <= a42[4];
					284:word <= a42[5];
					283:word <= a42[6];
					282:word <= a42[7];
					281:word <= a42[8];
					280:word <= a42[9];
					279:word <= a42[10];
					278:word <= a42[11];
					277:word <= a42[12];
					276:word <= a42[13];
					275:word <= a42[14];
					274:word <= a42[15];
					273:word <= a42[16];
					272:word <= a42[17];
					271:word <= a42[18];
					270:word <= a42[19];
					269:word <= a42[20];
					268:word <= a42[21];
					267:word <= a42[22];
					266:word <= a42[23];
					265:word <= a42[24];
					264:word <= a42[25];
					263:word <= a42[26];
					262:word <= a42[27];
					261:word <= a42[28];
					260:word <= a42[29];
					259:word <= a42[30];
					258:word <= a42[31];
					257:word <= a42[32];
					256:word <= a42[33];
					255:word <= a42[34];
					254:word <= a42[35];
					253:word <= a42[36];
					252:word <= a42[37];
					251:word <= a42[38];
					250:word <= a42[39];
					249:word <= a42[40];
					248:word <= a42[41];
					247:word <= a42[42];
					246:word <= a42[43];
					245:word <= a42[44];
					244:word <= a42[45];
					243:word <= a42[46];
					242:word <= a42[47];
					241:word <= a42[48];
					240:word <= a42[49];
					239:word <= a42[50];
					238:word <= a42[51];
					237:word <= a42[52];
					236:word <= a42[53];
					235:word <= a42[54];
					234:word <= a42[55];
					233:word <= a42[56];
					232:word <= a42[57];
					231:word <= a42[58];
					230:word <= a42[59];
					229:word <= a42[60];
					228:word <= a42[61];
					227:word <= a42[62];
					226:word <= a42[63];
					225:word <= a42[64];
					224:word <= a42[65];
					223:word <= a42[66];
					222:word <= a42[67];
					221:word <= a42[68];
					220:word <= a42[69];
					219:word <= a42[70];
					218:word <= a42[71];
					217:word <= a42[72];
					216:word <= a42[73];
					215:word <= a42[74];
					214:word <= a42[75];
					213:word <= a42[76];
					212:word <= a42[77];
					211:word <= a42[78];
					default:word <= a42[79];
					endcase
				end
				83:begin
				case(x)
					290:word <= a43[0];
					289:word <= a43[1];
					287:word <= a43[2];
					286:word <= a43[3];
					285:word <= a43[4];
					284:word <= a43[5];
					283:word <= a43[6];
					282:word <= a43[7];
					281:word <= a43[8];
					280:word <= a43[9];
					279:word <= a43[10];
					278:word <= a43[11];
					277:word <= a43[12];
					276:word <= a43[13];
					275:word <= a43[14];
					274:word <= a43[15];
					273:word <= a43[16];
					272:word <= a43[17];
					271:word <= a43[18];
					270:word <= a43[19];
					269:word <= a43[20];
					268:word <= a43[21];
					267:word <= a43[22];
					266:word <= a43[23];
					265:word <= a43[24];
					264:word <= a43[25];
					263:word <= a43[26];
					262:word <= a43[27];
					261:word <= a43[28];
					260:word <= a43[29];
					259:word <= a43[30];
					258:word <= a43[31];
					257:word <= a43[32];
					256:word <= a43[33];
					255:word <= a43[34];
					254:word <= a43[35];
					253:word <= a43[36];
					252:word <= a43[37];
					251:word <= a43[38];
					250:word <= a43[39];
					249:word <= a43[40];
					248:word <= a43[41];
					247:word <= a43[42];
					246:word <= a43[43];
					245:word <= a43[44];
					244:word <= a43[45];
					243:word <= a43[46];
					242:word <= a43[47];
					241:word <= a43[48];
					240:word <= a43[49];
					239:word <= a43[50];
					238:word <= a43[51];
					237:word <= a43[52];
					236:word <= a43[53];
					235:word <= a43[54];
					234:word <= a43[55];
					233:word <= a43[56];
					232:word <= a43[57];
					231:word <= a43[58];
					230:word <= a43[59];
					229:word <= a43[60];
					228:word <= a43[61];
					227:word <= a43[62];
					226:word <= a43[63];
					225:word <= a43[64];
					224:word <= a43[65];
					223:word <= a43[66];
					222:word <= a43[67];
					221:word <= a43[68];
					220:word <= a43[69];
					219:word <= a43[70];
					218:word <= a43[71];
					217:word <= a43[72];
					216:word <= a43[73];
					215:word <= a43[74];
					214:word <= a43[75];
					213:word <= a43[76];
					212:word <= a43[77];
					211:word <= a43[78];
					default:word <= a43[79];
					endcase
				end
				84:begin
				case(x)
					290:word <= a44[0];
					289:word <= a44[1];
					287:word <= a44[2];
					286:word <= a44[3];
					285:word <= a44[4];
					284:word <= a44[5];
					283:word <= a44[6];
					282:word <= a44[7];
					281:word <= a44[8];
					280:word <= a44[9];
					279:word <= a44[10];
					278:word <= a44[11];
					277:word <= a44[12];
					276:word <= a44[13];
					275:word <= a44[14];
					274:word <= a44[15];
					273:word <= a44[16];
					272:word <= a44[17];
					271:word <= a44[18];
					270:word <= a44[19];
					269:word <= a44[20];
					268:word <= a44[21];
					267:word <= a44[22];
					266:word <= a44[23];
					265:word <= a44[24];
					264:word <= a44[25];
					263:word <= a44[26];
					262:word <= a44[27];
					261:word <= a44[28];
					260:word <= a44[29];
					259:word <= a44[30];
					258:word <= a44[31];
					257:word <= a44[32];
					256:word <= a44[33];
					255:word <= a44[34];
					254:word <= a44[35];
					253:word <= a44[36];
					252:word <= a44[37];
					251:word <= a44[38];
					250:word <= a44[39];
					249:word <= a44[40];
					248:word <= a44[41];
					247:word <= a44[42];
					246:word <= a44[43];
					245:word <= a44[44];
					244:word <= a44[45];
					243:word <= a44[46];
					242:word <= a44[47];
					241:word <= a44[48];
					240:word <= a44[49];
					239:word <= a44[50];
					238:word <= a44[51];
					237:word <= a44[52];
					236:word <= a44[53];
					235:word <= a44[54];
					234:word <= a44[55];
					233:word <= a44[56];
					232:word <= a44[57];
					231:word <= a44[58];
					230:word <= a44[59];
					229:word <= a44[60];
					228:word <= a44[61];
					227:word <= a44[62];
					226:word <= a44[63];
					225:word <= a44[64];
					224:word <= a44[65];
					223:word <= a44[66];
					222:word <= a44[67];
					221:word <= a44[68];
					220:word <= a44[69];
					219:word <= a44[70];
					218:word <= a44[71];
					217:word <= a44[72];
					216:word <= a44[73];
					215:word <= a44[74];
					214:word <= a44[75];
					213:word <= a44[76];
					212:word <= a44[77];
					211:word <= a44[78];
					default:word <= a44[79];
					endcase
				end
				85:begin
				case(x)
					290:word <= a45[0];
					289:word <= a45[1];
					287:word <= a45[2];
					286:word <= a45[3];
					285:word <= a45[4];
					284:word <= a45[5];
					283:word <= a45[6];
					282:word <= a45[7];
					281:word <= a45[8];
					280:word <= a45[9];
					279:word <= a45[10];
					278:word <= a45[11];
					277:word <= a45[12];
					276:word <= a45[13];
					275:word <= a45[14];
					274:word <= a45[15];
					273:word <= a45[16];
					272:word <= a45[17];
					271:word <= a45[18];
					270:word <= a45[19];
					269:word <= a45[20];
					268:word <= a45[21];
					267:word <= a45[22];
					266:word <= a45[23];
					265:word <= a45[24];
					264:word <= a45[25];
					263:word <= a45[26];
					262:word <= a45[27];
					261:word <= a45[28];
					260:word <= a45[29];
					259:word <= a45[30];
					258:word <= a45[31];
					257:word <= a45[32];
					256:word <= a45[33];
					255:word <= a45[34];
					254:word <= a45[35];
					253:word <= a45[36];
					252:word <= a45[37];
					251:word <= a45[38];
					250:word <= a45[39];
					249:word <= a45[40];
					248:word <= a45[41];
					247:word <= a45[42];
					246:word <= a45[43];
					245:word <= a45[44];
					244:word <= a45[45];
					243:word <= a45[46];
					242:word <= a45[47];
					241:word <= a45[48];
					240:word <= a45[49];
					239:word <= a45[50];
					238:word <= a45[51];
					237:word <= a45[52];
					236:word <= a45[53];
					235:word <= a45[54];
					234:word <= a45[55];
					233:word <= a45[56];
					232:word <= a45[57];
					231:word <= a45[58];
					230:word <= a45[59];
					229:word <= a45[60];
					228:word <= a45[61];
					227:word <= a45[62];
					226:word <= a45[63];
					225:word <= a45[64];
					224:word <= a45[65];
					223:word <= a45[66];
					222:word <= a45[67];
					221:word <= a45[68];
					220:word <= a45[69];
					219:word <= a45[70];
					218:word <= a45[71];
					217:word <= a45[72];
					216:word <= a45[73];
					215:word <= a45[74];
					214:word <= a45[75];
					213:word <= a45[76];
					212:word <= a45[77];
					211:word <= a45[78];
					default:word <= a45[79];
					endcase
				end
				86:begin
				case(x)
					290:word <= a46[0];
					289:word <= a46[1];
					287:word <= a46[2];
					286:word <= a46[3];
					285:word <= a46[4];
					284:word <= a46[5];
					283:word <= a46[6];
					282:word <= a46[7];
					281:word <= a46[8];
					280:word <= a46[9];
					279:word <= a46[10];
					278:word <= a46[11];
					277:word <= a46[12];
					276:word <= a46[13];
					275:word <= a46[14];
					274:word <= a46[15];
					273:word <= a46[16];
					272:word <= a46[17];
					271:word <= a46[18];
					270:word <= a46[19];
					269:word <= a46[20];
					268:word <= a46[21];
					267:word <= a46[22];
					266:word <= a46[23];
					265:word <= a46[24];
					264:word <= a46[25];
					263:word <= a46[26];
					262:word <= a46[27];
					261:word <= a46[28];
					260:word <= a46[29];
					259:word <= a46[30];
					258:word <= a46[31];
					257:word <= a46[32];
					256:word <= a46[33];
					255:word <= a46[34];
					254:word <= a46[35];
					253:word <= a46[36];
					252:word <= a46[37];
					251:word <= a46[38];
					250:word <= a46[39];
					249:word <= a46[40];
					248:word <= a46[41];
					247:word <= a46[42];
					246:word <= a46[43];
					245:word <= a46[44];
					244:word <= a46[45];
					243:word <= a46[46];
					242:word <= a46[47];
					241:word <= a46[48];
					240:word <= a46[49];
					239:word <= a46[50];
					238:word <= a46[51];
					237:word <= a46[52];
					236:word <= a46[53];
					235:word <= a46[54];
					234:word <= a46[55];
					233:word <= a46[56];
					232:word <= a46[57];
					231:word <= a46[58];
					230:word <= a46[59];
					229:word <= a46[60];
					228:word <= a46[61];
					227:word <= a46[62];
					226:word <= a46[63];
					225:word <= a46[64];
					224:word <= a46[65];
					223:word <= a46[66];
					222:word <= a46[67];
					221:word <= a46[68];
					220:word <= a46[69];
					219:word <= a46[70];
					218:word <= a46[71];
					217:word <= a46[72];
					216:word <= a46[73];
					215:word <= a46[74];
					214:word <= a46[75];
					213:word <= a46[76];
					212:word <= a46[77];
					211:word <= a46[78];
					default:word <= a46[79];
					endcase
				end
				87:begin
				case(x)
					290:word <= a47[0];
					289:word <= a47[1];
					287:word <= a47[2];
					286:word <= a47[3];
					285:word <= a47[4];
					284:word <= a47[5];
					283:word <= a47[6];
					282:word <= a47[7];
					281:word <= a47[8];
					280:word <= a47[9];
					279:word <= a47[10];
					278:word <= a47[11];
					277:word <= a47[12];
					276:word <= a47[13];
					275:word <= a47[14];
					274:word <= a47[15];
					273:word <= a47[16];
					272:word <= a47[17];
					271:word <= a47[18];
					270:word <= a47[19];
					269:word <= a47[20];
					268:word <= a47[21];
					267:word <= a47[22];
					266:word <= a47[23];
					265:word <= a47[24];
					264:word <= a47[25];
					263:word <= a47[26];
					262:word <= a47[27];
					261:word <= a47[28];
					260:word <= a47[29];
					259:word <= a47[30];
					258:word <= a47[31];
					257:word <= a47[32];
					256:word <= a47[33];
					255:word <= a47[34];
					254:word <= a47[35];
					253:word <= a47[36];
					252:word <= a47[37];
					251:word <= a47[38];
					250:word <= a47[39];
					249:word <= a47[40];
					248:word <= a47[41];
					247:word <= a47[42];
					246:word <= a47[43];
					245:word <= a47[44];
					244:word <= a47[45];
					243:word <= a47[46];
					242:word <= a47[47];
					241:word <= a47[48];
					240:word <= a47[49];
					239:word <= a47[50];
					238:word <= a47[51];
					237:word <= a47[52];
					236:word <= a47[53];
					235:word <= a47[54];
					234:word <= a47[55];
					233:word <= a47[56];
					232:word <= a47[57];
					231:word <= a47[58];
					230:word <= a47[59];
					229:word <= a47[60];
					228:word <= a47[61];
					227:word <= a47[62];
					226:word <= a47[63];
					225:word <= a47[64];
					224:word <= a47[65];
					223:word <= a47[66];
					222:word <= a47[67];
					221:word <= a47[68];
					220:word <= a47[69];
					219:word <= a47[70];
					218:word <= a47[71];
					217:word <= a47[72];
					216:word <= a47[73];
					215:word <= a47[74];
					214:word <= a47[75];
					213:word <= a47[76];
					212:word <= a47[77];
					211:word <= a47[78];
					default:word <= a47[79];
					endcase
				end
				88:begin
				case(x)
					290:word <= a48[0];
					289:word <= a48[1];
					287:word <= a48[2];
					286:word <= a48[3];
					285:word <= a48[4];
					284:word <= a48[5];
					283:word <= a48[6];
					282:word <= a48[7];
					281:word <= a48[8];
					280:word <= a48[9];
					279:word <= a48[10];
					278:word <= a48[11];
					277:word <= a48[12];
					276:word <= a48[13];
					275:word <= a48[14];
					274:word <= a48[15];
					273:word <= a48[16];
					272:word <= a48[17];
					271:word <= a48[18];
					270:word <= a48[19];
					269:word <= a48[20];
					268:word <= a48[21];
					267:word <= a48[22];
					266:word <= a48[23];
					265:word <= a48[24];
					264:word <= a48[25];
					263:word <= a48[26];
					262:word <= a48[27];
					261:word <= a48[28];
					260:word <= a48[29];
					259:word <= a48[30];
					258:word <= a48[31];
					257:word <= a48[32];
					256:word <= a48[33];
					255:word <= a48[34];
					254:word <= a48[35];
					253:word <= a48[36];
					252:word <= a48[37];
					251:word <= a48[38];
					250:word <= a48[39];
					249:word <= a48[40];
					248:word <= a48[41];
					247:word <= a48[42];
					246:word <= a48[43];
					245:word <= a48[44];
					244:word <= a48[45];
					243:word <= a48[46];
					242:word <= a48[47];
					241:word <= a48[48];
					240:word <= a48[49];
					239:word <= a48[50];
					238:word <= a48[51];
					237:word <= a48[52];
					236:word <= a48[53];
					235:word <= a48[54];
					234:word <= a48[55];
					233:word <= a48[56];
					232:word <= a48[57];
					231:word <= a48[58];
					230:word <= a48[59];
					229:word <= a48[60];
					228:word <= a48[61];
					227:word <= a48[62];
					226:word <= a48[63];
					225:word <= a48[64];
					224:word <= a48[65];
					223:word <= a48[66];
					222:word <= a48[67];
					221:word <= a48[68];
					220:word <= a48[69];
					219:word <= a48[70];
					218:word <= a48[71];
					217:word <= a48[72];
					216:word <= a48[73];
					215:word <= a48[74];
					214:word <= a48[75];
					213:word <= a48[76];
					212:word <= a48[77];
					211:word <= a48[78];
					default:word <= a48[79];
					endcase
				end
				89:begin
				case(x)
					290:word <= a49[0];
					289:word <= a49[1];
					287:word <= a49[2];
					286:word <= a49[3];
					285:word <= a49[4];
					284:word <= a49[5];
					283:word <= a49[6];
					282:word <= a49[7];
					281:word <= a49[8];
					280:word <= a49[9];
					279:word <= a49[10];
					278:word <= a49[11];
					277:word <= a49[12];
					276:word <= a49[13];
					275:word <= a49[14];
					274:word <= a49[15];
					273:word <= a49[16];
					272:word <= a49[17];
					271:word <= a49[18];
					270:word <= a49[19];
					269:word <= a49[20];
					268:word <= a49[21];
					267:word <= a49[22];
					266:word <= a49[23];
					265:word <= a49[24];
					264:word <= a49[25];
					263:word <= a49[26];
					262:word <= a49[27];
					261:word <= a49[28];
					260:word <= a49[29];
					259:word <= a49[30];
					258:word <= a49[31];
					257:word <= a49[32];
					256:word <= a49[33];
					255:word <= a49[34];
					254:word <= a49[35];
					253:word <= a49[36];
					252:word <= a49[37];
					251:word <= a49[38];
					250:word <= a49[39];
					249:word <= a49[40];
					248:word <= a49[41];
					247:word <= a49[42];
					246:word <= a49[43];
					245:word <= a49[44];
					244:word <= a49[45];
					243:word <= a49[46];
					242:word <= a49[47];
					241:word <= a49[48];
					240:word <= a49[49];
					239:word <= a49[50];
					238:word <= a49[51];
					237:word <= a49[52];
					236:word <= a49[53];
					235:word <= a49[54];
					234:word <= a49[55];
					233:word <= a49[56];
					232:word <= a49[57];
					231:word <= a49[58];
					230:word <= a49[59];
					229:word <= a49[60];
					228:word <= a49[61];
					227:word <= a49[62];
					226:word <= a49[63];
					225:word <= a49[64];
					224:word <= a49[65];
					223:word <= a49[66];
					222:word <= a49[67];
					221:word <= a49[68];
					220:word <= a49[69];
					219:word <= a49[70];
					218:word <= a49[71];
					217:word <= a49[72];
					216:word <= a49[73];
					215:word <= a49[74];
					214:word <= a49[75];
					213:word <= a49[76];
					212:word <= a49[77];
					211:word <= a49[78];
					default:word <= a49[79];
					endcase
				end
				90:begin
				case(x)
					290:word <= a50[0];
					289:word <= a50[1];
					287:word <= a50[2];
					286:word <= a50[3];
					285:word <= a50[4];
					284:word <= a50[5];
					283:word <= a50[6];
					282:word <= a50[7];
					281:word <= a50[8];
					280:word <= a50[9];
					279:word <= a50[10];
					278:word <= a50[11];
					277:word <= a50[12];
					276:word <= a50[13];
					275:word <= a50[14];
					274:word <= a50[15];
					273:word <= a50[16];
					272:word <= a50[17];
					271:word <= a50[18];
					270:word <= a50[19];
					269:word <= a50[20];
					268:word <= a50[21];
					267:word <= a50[22];
					266:word <= a50[23];
					265:word <= a50[24];
					264:word <= a50[25];
					263:word <= a50[26];
					262:word <= a50[27];
					261:word <= a50[28];
					260:word <= a50[29];
					259:word <= a50[30];
					258:word <= a50[31];
					257:word <= a50[32];
					256:word <= a50[33];
					255:word <= a50[34];
					254:word <= a50[35];
					253:word <= a50[36];
					252:word <= a50[37];
					251:word <= a50[38];
					250:word <= a50[39];
					249:word <= a50[40];
					248:word <= a50[41];
					247:word <= a50[42];
					246:word <= a50[43];
					245:word <= a50[44];
					244:word <= a50[45];
					243:word <= a50[46];
					242:word <= a50[47];
					241:word <= a50[48];
					240:word <= a50[49];
					239:word <= a50[50];
					238:word <= a50[51];
					237:word <= a50[52];
					236:word <= a50[53];
					235:word <= a50[54];
					234:word <= a50[55];
					233:word <= a50[56];
					232:word <= a50[57];
					231:word <= a50[58];
					230:word <= a50[59];
					229:word <= a50[60];
					228:word <= a50[61];
					227:word <= a50[62];
					226:word <= a50[63];
					225:word <= a50[64];
					224:word <= a50[65];
					223:word <= a50[66];
					222:word <= a50[67];
					221:word <= a50[68];
					220:word <= a50[69];
					219:word <= a50[70];
					218:word <= a50[71];
					217:word <= a50[72];
					216:word <= a50[73];
					215:word <= a50[74];
					214:word <= a50[75];
					213:word <= a50[76];
					212:word <= a50[77];
					211:word <= a50[78];
					default:word <= a50[79];
					endcase
				end
				91:begin
				case(x)
					290:word <= a51[0];
					289:word <= a51[1];
					287:word <= a51[2];
					286:word <= a51[3];
					285:word <= a51[4];
					284:word <= a51[5];
					283:word <= a51[6];
					282:word <= a51[7];
					281:word <= a51[8];
					280:word <= a51[9];
					279:word <= a51[10];
					278:word <= a51[11];
					277:word <= a51[12];
					276:word <= a51[13];
					275:word <= a51[14];
					274:word <= a51[15];
					273:word <= a51[16];
					272:word <= a51[17];
					271:word <= a51[18];
					270:word <= a51[19];
					269:word <= a51[20];
					268:word <= a51[21];
					267:word <= a51[22];
					266:word <= a51[23];
					265:word <= a51[24];
					264:word <= a51[25];
					263:word <= a51[26];
					262:word <= a51[27];
					261:word <= a51[28];
					260:word <= a51[29];
					259:word <= a51[30];
					258:word <= a51[31];
					257:word <= a51[32];
					256:word <= a51[33];
					255:word <= a51[34];
					254:word <= a51[35];
					253:word <= a51[36];
					252:word <= a51[37];
					251:word <= a51[38];
					250:word <= a51[39];
					249:word <= a51[40];
					248:word <= a51[41];
					247:word <= a51[42];
					246:word <= a51[43];
					245:word <= a51[44];
					244:word <= a51[45];
					243:word <= a51[46];
					242:word <= a51[47];
					241:word <= a51[48];
					240:word <= a51[49];
					239:word <= a51[50];
					238:word <= a51[51];
					237:word <= a51[52];
					236:word <= a51[53];
					235:word <= a51[54];
					234:word <= a51[55];
					233:word <= a51[56];
					232:word <= a51[57];
					231:word <= a51[58];
					230:word <= a51[59];
					229:word <= a51[60];
					228:word <= a51[61];
					227:word <= a51[62];
					226:word <= a51[63];
					225:word <= a51[64];
					224:word <= a51[65];
					223:word <= a51[66];
					222:word <= a51[67];
					221:word <= a51[68];
					220:word <= a51[69];
					219:word <= a51[70];
					218:word <= a51[71];
					217:word <= a51[72];
					216:word <= a51[73];
					215:word <= a51[74];
					214:word <= a51[75];
					213:word <= a51[76];
					212:word <= a51[77];
					211:word <= a51[78];
					default:word <= a51[79];
					endcase
				end
				92:begin
				case(x)
					290:word <= a52[0];
					289:word <= a52[1];
					287:word <= a52[2];
					286:word <= a52[3];
					285:word <= a52[4];
					284:word <= a52[5];
					283:word <= a52[6];
					282:word <= a52[7];
					281:word <= a52[8];
					280:word <= a52[9];
					279:word <= a52[10];
					278:word <= a52[11];
					277:word <= a52[12];
					276:word <= a52[13];
					275:word <= a52[14];
					274:word <= a52[15];
					273:word <= a52[16];
					272:word <= a52[17];
					271:word <= a52[18];
					270:word <= a52[19];
					269:word <= a52[20];
					268:word <= a52[21];
					267:word <= a52[22];
					266:word <= a52[23];
					265:word <= a52[24];
					264:word <= a52[25];
					263:word <= a52[26];
					262:word <= a52[27];
					261:word <= a52[28];
					260:word <= a52[29];
					259:word <= a52[30];
					258:word <= a52[31];
					257:word <= a52[32];
					256:word <= a52[33];
					255:word <= a52[34];
					254:word <= a52[35];
					253:word <= a52[36];
					252:word <= a52[37];
					251:word <= a52[38];
					250:word <= a52[39];
					249:word <= a52[40];
					248:word <= a52[41];
					247:word <= a52[42];
					246:word <= a52[43];
					245:word <= a52[44];
					244:word <= a52[45];
					243:word <= a52[46];
					242:word <= a52[47];
					241:word <= a52[48];
					240:word <= a52[49];
					239:word <= a52[50];
					238:word <= a52[51];
					237:word <= a52[52];
					236:word <= a52[53];
					235:word <= a52[54];
					234:word <= a52[55];
					233:word <= a52[56];
					232:word <= a52[57];
					231:word <= a52[58];
					230:word <= a52[59];
					229:word <= a52[60];
					228:word <= a52[61];
					227:word <= a52[62];
					226:word <= a52[63];
					225:word <= a52[64];
					224:word <= a52[65];
					223:word <= a52[66];
					222:word <= a52[67];
					221:word <= a52[68];
					220:word <= a52[69];
					219:word <= a52[70];
					218:word <= a52[71];
					217:word <= a52[72];
					216:word <= a52[73];
					215:word <= a52[74];
					214:word <= a52[75];
					213:word <= a52[76];
					212:word <= a52[77];
					211:word <= a52[78];
					default:word <= a52[79];
					endcase
				end
				93:begin
				case(x)
					290:word <= a53[0];
					289:word <= a53[1];
					287:word <= a53[2];
					286:word <= a53[3];
					285:word <= a53[4];
					284:word <= a53[5];
					283:word <= a53[6];
					282:word <= a53[7];
					281:word <= a53[8];
					280:word <= a53[9];
					279:word <= a53[10];
					278:word <= a53[11];
					277:word <= a53[12];
					276:word <= a53[13];
					275:word <= a53[14];
					274:word <= a53[15];
					273:word <= a53[16];
					272:word <= a53[17];
					271:word <= a53[18];
					270:word <= a53[19];
					269:word <= a53[20];
					268:word <= a53[21];
					267:word <= a53[22];
					266:word <= a53[23];
					265:word <= a53[24];
					264:word <= a53[25];
					263:word <= a53[26];
					262:word <= a53[27];
					261:word <= a53[28];
					260:word <= a53[29];
					259:word <= a53[30];
					258:word <= a53[31];
					257:word <= a53[32];
					256:word <= a53[33];
					255:word <= a53[34];
					254:word <= a53[35];
					253:word <= a53[36];
					252:word <= a53[37];
					251:word <= a53[38];
					250:word <= a53[39];
					249:word <= a53[40];
					248:word <= a53[41];
					247:word <= a53[42];
					246:word <= a53[43];
					245:word <= a53[44];
					244:word <= a53[45];
					243:word <= a53[46];
					242:word <= a53[47];
					241:word <= a53[48];
					240:word <= a53[49];
					239:word <= a53[50];
					238:word <= a53[51];
					237:word <= a53[52];
					236:word <= a53[53];
					235:word <= a53[54];
					234:word <= a53[55];
					233:word <= a53[56];
					232:word <= a53[57];
					231:word <= a53[58];
					230:word <= a53[59];
					229:word <= a53[60];
					228:word <= a53[61];
					227:word <= a53[62];
					226:word <= a53[63];
					225:word <= a53[64];
					224:word <= a53[65];
					223:word <= a53[66];
					222:word <= a53[67];
					221:word <= a53[68];
					220:word <= a53[69];
					219:word <= a53[70];
					218:word <= a53[71];
					217:word <= a53[72];
					216:word <= a53[73];
					215:word <= a53[74];
					214:word <= a53[75];
					213:word <= a53[76];
					212:word <= a53[77];
					211:word <= a53[78];
					default:word <= a53[79];
					endcase
				end
				94:begin
				case(x)
					290:word <= a54[0];
					289:word <= a54[1];
					287:word <= a54[2];
					286:word <= a54[3];
					285:word <= a54[4];
					284:word <= a54[5];
					283:word <= a54[6];
					282:word <= a54[7];
					281:word <= a54[8];
					280:word <= a54[9];
					279:word <= a54[10];
					278:word <= a54[11];
					277:word <= a54[12];
					276:word <= a54[13];
					275:word <= a54[14];
					274:word <= a54[15];
					273:word <= a54[16];
					272:word <= a54[17];
					271:word <= a54[18];
					270:word <= a54[19];
					269:word <= a54[20];
					268:word <= a54[21];
					267:word <= a54[22];
					266:word <= a54[23];
					265:word <= a54[24];
					264:word <= a54[25];
					263:word <= a54[26];
					262:word <= a54[27];
					261:word <= a54[28];
					260:word <= a54[29];
					259:word <= a54[30];
					258:word <= a54[31];
					257:word <= a54[32];
					256:word <= a54[33];
					255:word <= a54[34];
					254:word <= a54[35];
					253:word <= a54[36];
					252:word <= a54[37];
					251:word <= a54[38];
					250:word <= a54[39];
					249:word <= a54[40];
					248:word <= a54[41];
					247:word <= a54[42];
					246:word <= a54[43];
					245:word <= a54[44];
					244:word <= a54[45];
					243:word <= a54[46];
					242:word <= a54[47];
					241:word <= a54[48];
					240:word <= a54[49];
					239:word <= a54[50];
					238:word <= a54[51];
					237:word <= a54[52];
					236:word <= a54[53];
					235:word <= a54[54];
					234:word <= a54[55];
					233:word <= a54[56];
					232:word <= a54[57];
					231:word <= a54[58];
					230:word <= a54[59];
					229:word <= a54[60];
					228:word <= a54[61];
					227:word <= a54[62];
					226:word <= a54[63];
					225:word <= a54[64];
					224:word <= a54[65];
					223:word <= a54[66];
					222:word <= a54[67];
					221:word <= a54[68];
					220:word <= a54[69];
					219:word <= a54[70];
					218:word <= a54[71];
					217:word <= a54[72];
					216:word <= a54[73];
					215:word <= a54[74];
					214:word <= a54[75];
					213:word <= a54[76];
					212:word <= a54[77];
					211:word <= a54[78];
					default:word <= a54[79];
					endcase
				end
				95:begin
				case(x)
					290:word <= a55[0];
					289:word <= a55[1];
					287:word <= a55[2];
					286:word <= a55[3];
					285:word <= a55[4];
					284:word <= a55[5];
					283:word <= a55[6];
					282:word <= a55[7];
					281:word <= a55[8];
					280:word <= a55[9];
					279:word <= a55[10];
					278:word <= a55[11];
					277:word <= a55[12];
					276:word <= a55[13];
					275:word <= a55[14];
					274:word <= a55[15];
					273:word <= a55[16];
					272:word <= a55[17];
					271:word <= a55[18];
					270:word <= a55[19];
					269:word <= a55[20];
					268:word <= a55[21];
					267:word <= a55[22];
					266:word <= a55[23];
					265:word <= a55[24];
					264:word <= a55[25];
					263:word <= a55[26];
					262:word <= a55[27];
					261:word <= a55[28];
					260:word <= a55[29];
					259:word <= a55[30];
					258:word <= a55[31];
					257:word <= a55[32];
					256:word <= a55[33];
					255:word <= a55[34];
					254:word <= a55[35];
					253:word <= a55[36];
					252:word <= a55[37];
					251:word <= a55[38];
					250:word <= a55[39];
					249:word <= a55[40];
					248:word <= a55[41];
					247:word <= a55[42];
					246:word <= a55[43];
					245:word <= a55[44];
					244:word <= a55[45];
					243:word <= a55[46];
					242:word <= a55[47];
					241:word <= a55[48];
					240:word <= a55[49];
					239:word <= a55[50];
					238:word <= a55[51];
					237:word <= a55[52];
					236:word <= a55[53];
					235:word <= a55[54];
					234:word <= a55[55];
					233:word <= a55[56];
					232:word <= a55[57];
					231:word <= a55[58];
					230:word <= a55[59];
					229:word <= a55[60];
					228:word <= a55[61];
					227:word <= a55[62];
					226:word <= a55[63];
					225:word <= a55[64];
					224:word <= a55[65];
					223:word <= a55[66];
					222:word <= a55[67];
					221:word <= a55[68];
					220:word <= a55[69];
					219:word <= a55[70];
					218:word <= a55[71];
					217:word <= a55[72];
					216:word <= a55[73];
					215:word <= a55[74];
					214:word <= a55[75];
					213:word <= a55[76];
					212:word <= a55[77];
					211:word <= a55[78];
					default:word <= a55[79];
					endcase
				end
				96:begin
				case(x)
					290:word <= a56[0];
					289:word <= a56[1];
					287:word <= a56[2];
					286:word <= a56[3];
					285:word <= a56[4];
					284:word <= a56[5];
					283:word <= a56[6];
					282:word <= a56[7];
					281:word <= a56[8];
					280:word <= a56[9];
					279:word <= a56[10];
					278:word <= a56[11];
					277:word <= a56[12];
					276:word <= a56[13];
					275:word <= a56[14];
					274:word <= a56[15];
					273:word <= a56[16];
					272:word <= a56[17];
					271:word <= a56[18];
					270:word <= a56[19];
					269:word <= a56[20];
					268:word <= a56[21];
					267:word <= a56[22];
					266:word <= a56[23];
					265:word <= a56[24];
					264:word <= a56[25];
					263:word <= a56[26];
					262:word <= a56[27];
					261:word <= a56[28];
					260:word <= a56[29];
					259:word <= a56[30];
					258:word <= a56[31];
					257:word <= a56[32];
					256:word <= a56[33];
					255:word <= a56[34];
					254:word <= a56[35];
					253:word <= a56[36];
					252:word <= a56[37];
					251:word <= a56[38];
					250:word <= a56[39];
					249:word <= a56[40];
					248:word <= a56[41];
					247:word <= a56[42];
					246:word <= a56[43];
					245:word <= a56[44];
					244:word <= a56[45];
					243:word <= a56[46];
					242:word <= a56[47];
					241:word <= a56[48];
					240:word <= a56[49];
					239:word <= a56[50];
					238:word <= a56[51];
					237:word <= a56[52];
					236:word <= a56[53];
					235:word <= a56[54];
					234:word <= a56[55];
					233:word <= a56[56];
					232:word <= a56[57];
					231:word <= a56[58];
					230:word <= a56[59];
					229:word <= a56[60];
					228:word <= a56[61];
					227:word <= a56[62];
					226:word <= a56[63];
					225:word <= a56[64];
					224:word <= a56[65];
					223:word <= a56[66];
					222:word <= a56[67];
					221:word <= a56[68];
					220:word <= a56[69];
					219:word <= a56[70];
					218:word <= a56[71];
					217:word <= a56[72];
					216:word <= a56[73];
					215:word <= a56[74];
					214:word <= a56[75];
					213:word <= a56[76];
					212:word <= a56[77];
					211:word <= a56[78];
					default:word <= a56[79];
					endcase
				end
				97:begin
				case(x)
					290:word <= a57[0];
					289:word <= a57[1];
					287:word <= a57[2];
					286:word <= a57[3];
					285:word <= a57[4];
					284:word <= a57[5];
					283:word <= a57[6];
					282:word <= a57[7];
					281:word <= a57[8];
					280:word <= a57[9];
					279:word <= a57[10];
					278:word <= a57[11];
					277:word <= a57[12];
					276:word <= a57[13];
					275:word <= a57[14];
					274:word <= a57[15];
					273:word <= a57[16];
					272:word <= a57[17];
					271:word <= a57[18];
					270:word <= a57[19];
					269:word <= a57[20];
					268:word <= a57[21];
					267:word <= a57[22];
					266:word <= a57[23];
					265:word <= a57[24];
					264:word <= a57[25];
					263:word <= a57[26];
					262:word <= a57[27];
					261:word <= a57[28];
					260:word <= a57[29];
					259:word <= a57[30];
					258:word <= a57[31];
					257:word <= a57[32];
					256:word <= a57[33];
					255:word <= a57[34];
					254:word <= a57[35];
					253:word <= a57[36];
					252:word <= a57[37];
					251:word <= a57[38];
					250:word <= a57[39];
					249:word <= a57[40];
					248:word <= a57[41];
					247:word <= a57[42];
					246:word <= a57[43];
					245:word <= a57[44];
					244:word <= a57[45];
					243:word <= a57[46];
					242:word <= a57[47];
					241:word <= a57[48];
					240:word <= a57[49];
					239:word <= a57[50];
					238:word <= a57[51];
					237:word <= a57[52];
					236:word <= a57[53];
					235:word <= a57[54];
					234:word <= a57[55];
					233:word <= a57[56];
					232:word <= a57[57];
					231:word <= a57[58];
					230:word <= a57[59];
					229:word <= a57[60];
					228:word <= a57[61];
					227:word <= a57[62];
					226:word <= a57[63];
					225:word <= a57[64];
					224:word <= a57[65];
					223:word <= a57[66];
					222:word <= a57[67];
					221:word <= a57[68];
					220:word <= a57[69];
					219:word <= a57[70];
					218:word <= a57[71];
					217:word <= a57[72];
					216:word <= a57[73];
					215:word <= a57[74];
					214:word <= a57[75];
					213:word <= a57[76];
					212:word <= a57[77];
					211:word <= a57[78];
					default:word <= a57[79];
					endcase
				end
				98:begin
				case(x)
					290:word <= a58[0];
					289:word <= a58[1];
					287:word <= a58[2];
					286:word <= a58[3];
					285:word <= a58[4];
					284:word <= a58[5];
					283:word <= a58[6];
					282:word <= a58[7];
					281:word <= a58[8];
					280:word <= a58[9];
					279:word <= a58[10];
					278:word <= a58[11];
					277:word <= a58[12];
					276:word <= a58[13];
					275:word <= a58[14];
					274:word <= a58[15];
					273:word <= a58[16];
					272:word <= a58[17];
					271:word <= a58[18];
					270:word <= a58[19];
					269:word <= a58[20];
					268:word <= a58[21];
					267:word <= a58[22];
					266:word <= a58[23];
					265:word <= a58[24];
					264:word <= a58[25];
					263:word <= a58[26];
					262:word <= a58[27];
					261:word <= a58[28];
					260:word <= a58[29];
					259:word <= a58[30];
					258:word <= a58[31];
					257:word <= a58[32];
					256:word <= a58[33];
					255:word <= a58[34];
					254:word <= a58[35];
					253:word <= a58[36];
					252:word <= a58[37];
					251:word <= a58[38];
					250:word <= a58[39];
					249:word <= a58[40];
					248:word <= a58[41];
					247:word <= a58[42];
					246:word <= a58[43];
					245:word <= a58[44];
					244:word <= a58[45];
					243:word <= a58[46];
					242:word <= a58[47];
					241:word <= a58[48];
					240:word <= a58[49];
					239:word <= a58[50];
					238:word <= a58[51];
					237:word <= a58[52];
					236:word <= a58[53];
					235:word <= a58[54];
					234:word <= a58[55];
					233:word <= a58[56];
					232:word <= a58[57];
					231:word <= a58[58];
					230:word <= a58[59];
					229:word <= a58[60];
					228:word <= a58[61];
					227:word <= a58[62];
					226:word <= a58[63];
					225:word <= a58[64];
					224:word <= a58[65];
					223:word <= a58[66];
					222:word <= a58[67];
					221:word <= a58[68];
					220:word <= a58[69];
					219:word <= a58[70];
					218:word <= a58[71];
					217:word <= a58[72];
					216:word <= a58[73];
					215:word <= a58[74];
					214:word <= a58[75];
					213:word <= a58[76];
					212:word <= a58[77];
					211:word <= a58[78];
					default:word <= a58[79];
					endcase
				end
				99:begin
				case(x)
					290:word <= a59[0];
					289:word <= a59[1];
					287:word <= a59[2];
					286:word <= a59[3];
					285:word <= a59[4];
					284:word <= a59[5];
					283:word <= a59[6];
					282:word <= a59[7];
					281:word <= a59[8];
					280:word <= a59[9];
					279:word <= a59[10];
					278:word <= a59[11];
					277:word <= a59[12];
					276:word <= a59[13];
					275:word <= a59[14];
					274:word <= a59[15];
					273:word <= a59[16];
					272:word <= a59[17];
					271:word <= a59[18];
					270:word <= a59[19];
					269:word <= a59[20];
					268:word <= a59[21];
					267:word <= a59[22];
					266:word <= a59[23];
					265:word <= a59[24];
					264:word <= a59[25];
					263:word <= a59[26];
					262:word <= a59[27];
					261:word <= a59[28];
					260:word <= a59[29];
					259:word <= a59[30];
					258:word <= a59[31];
					257:word <= a59[32];
					256:word <= a59[33];
					255:word <= a59[34];
					254:word <= a59[35];
					253:word <= a59[36];
					252:word <= a59[37];
					251:word <= a59[38];
					250:word <= a59[39];
					249:word <= a59[40];
					248:word <= a59[41];
					247:word <= a59[42];
					246:word <= a59[43];
					245:word <= a59[44];
					244:word <= a59[45];
					243:word <= a59[46];
					242:word <= a59[47];
					241:word <= a59[48];
					240:word <= a59[49];
					239:word <= a59[50];
					238:word <= a59[51];
					237:word <= a59[52];
					236:word <= a59[53];
					235:word <= a59[54];
					234:word <= a59[55];
					233:word <= a59[56];
					232:word <= a59[57];
					231:word <= a59[58];
					230:word <= a59[59];
					229:word <= a59[60];
					228:word <= a59[61];
					227:word <= a59[62];
					226:word <= a59[63];
					225:word <= a59[64];
					224:word <= a59[65];
					223:word <= a59[66];
					222:word <= a59[67];
					221:word <= a59[68];
					220:word <= a59[69];
					219:word <= a59[70];
					218:word <= a59[71];
					217:word <= a59[72];
					216:word <= a59[73];
					215:word <= a59[74];
					214:word <= a59[75];
					213:word <= a59[76];
					212:word <= a59[77];
					211:word <= a59[78];
					default:word <= a59[79];
					endcase
				end
				100:begin
				case(x)
					290:word <= a60[0];
					289:word <= a60[1];
					287:word <= a60[2];
					286:word <= a60[3];
					285:word <= a60[4];
					284:word <= a60[5];
					283:word <= a60[6];
					282:word <= a60[7];
					281:word <= a60[8];
					280:word <= a60[9];
					279:word <= a60[10];
					278:word <= a60[11];
					277:word <= a60[12];
					276:word <= a60[13];
					275:word <= a60[14];
					274:word <= a60[15];
					273:word <= a60[16];
					272:word <= a60[17];
					271:word <= a60[18];
					270:word <= a60[19];
					269:word <= a60[20];
					268:word <= a60[21];
					267:word <= a60[22];
					266:word <= a60[23];
					265:word <= a60[24];
					264:word <= a60[25];
					263:word <= a60[26];
					262:word <= a60[27];
					261:word <= a60[28];
					260:word <= a60[29];
					259:word <= a60[30];
					258:word <= a60[31];
					257:word <= a60[32];
					256:word <= a60[33];
					255:word <= a60[34];
					254:word <= a60[35];
					253:word <= a60[36];
					252:word <= a60[37];
					251:word <= a60[38];
					250:word <= a60[39];
					249:word <= a60[40];
					248:word <= a60[41];
					247:word <= a60[42];
					246:word <= a60[43];
					245:word <= a60[44];
					244:word <= a60[45];
					243:word <= a60[46];
					242:word <= a60[47];
					241:word <= a60[48];
					240:word <= a60[49];
					239:word <= a60[50];
					238:word <= a60[51];
					237:word <= a60[52];
					236:word <= a60[53];
					235:word <= a60[54];
					234:word <= a60[55];
					233:word <= a60[56];
					232:word <= a60[57];
					231:word <= a60[58];
					230:word <= a60[59];
					229:word <= a60[60];
					228:word <= a60[61];
					227:word <= a60[62];
					226:word <= a60[63];
					225:word <= a60[64];
					224:word <= a60[65];
					223:word <= a60[66];
					222:word <= a60[67];
					221:word <= a60[68];
					220:word <= a60[69];
					219:word <= a60[70];
					218:word <= a60[71];
					217:word <= a60[72];
					216:word <= a60[73];
					215:word <= a60[74];
					214:word <= a60[75];
					213:word <= a60[76];
					212:word <= a60[77];
					211:word <= a60[78];
					default:word <= a60[79];
					endcase
				end
				101:begin
				case(x)
					290:word <= a61[0];
					289:word <= a61[1];
					287:word <= a61[2];
					286:word <= a61[3];
					285:word <= a61[4];
					284:word <= a61[5];
					283:word <= a61[6];
					282:word <= a61[7];
					281:word <= a61[8];
					280:word <= a61[9];
					279:word <= a61[10];
					278:word <= a61[11];
					277:word <= a61[12];
					276:word <= a61[13];
					275:word <= a61[14];
					274:word <= a61[15];
					273:word <= a61[16];
					272:word <= a61[17];
					271:word <= a61[18];
					270:word <= a61[19];
					269:word <= a61[20];
					268:word <= a61[21];
					267:word <= a61[22];
					266:word <= a61[23];
					265:word <= a61[24];
					264:word <= a61[25];
					263:word <= a61[26];
					262:word <= a61[27];
					261:word <= a61[28];
					260:word <= a61[29];
					259:word <= a61[30];
					258:word <= a61[31];
					257:word <= a61[32];
					256:word <= a61[33];
					255:word <= a61[34];
					254:word <= a61[35];
					253:word <= a61[36];
					252:word <= a61[37];
					251:word <= a61[38];
					250:word <= a61[39];
					249:word <= a61[40];
					248:word <= a61[41];
					247:word <= a61[42];
					246:word <= a61[43];
					245:word <= a61[44];
					244:word <= a61[45];
					243:word <= a61[46];
					242:word <= a61[47];
					241:word <= a61[48];
					240:word <= a61[49];
					239:word <= a61[50];
					238:word <= a61[51];
					237:word <= a61[52];
					236:word <= a61[53];
					235:word <= a61[54];
					234:word <= a61[55];
					233:word <= a61[56];
					232:word <= a61[57];
					231:word <= a61[58];
					230:word <= a61[59];
					229:word <= a61[60];
					228:word <= a61[61];
					227:word <= a61[62];
					226:word <= a61[63];
					225:word <= a61[64];
					224:word <= a61[65];
					223:word <= a61[66];
					222:word <= a61[67];
					221:word <= a61[68];
					220:word <= a61[69];
					219:word <= a61[70];
					218:word <= a61[71];
					217:word <= a61[72];
					216:word <= a61[73];
					215:word <= a61[74];
					214:word <= a61[75];
					213:word <= a61[76];
					212:word <= a61[77];
					211:word <= a61[78];
					default:word <= a61[79];
					endcase
				end
				102:begin
				case(x)
					290:word <= a62[0];
					289:word <= a62[1];
					287:word <= a62[2];
					286:word <= a62[3];
					285:word <= a62[4];
					284:word <= a62[5];
					283:word <= a62[6];
					282:word <= a62[7];
					281:word <= a62[8];
					280:word <= a62[9];
					279:word <= a62[10];
					278:word <= a62[11];
					277:word <= a62[12];
					276:word <= a62[13];
					275:word <= a62[14];
					274:word <= a62[15];
					273:word <= a62[16];
					272:word <= a62[17];
					271:word <= a62[18];
					270:word <= a62[19];
					269:word <= a62[20];
					268:word <= a62[21];
					267:word <= a62[22];
					266:word <= a62[23];
					265:word <= a62[24];
					264:word <= a62[25];
					263:word <= a62[26];
					262:word <= a62[27];
					261:word <= a62[28];
					260:word <= a62[29];
					259:word <= a62[30];
					258:word <= a62[31];
					257:word <= a62[32];
					256:word <= a62[33];
					255:word <= a62[34];
					254:word <= a62[35];
					253:word <= a62[36];
					252:word <= a62[37];
					251:word <= a62[38];
					250:word <= a62[39];
					249:word <= a62[40];
					248:word <= a62[41];
					247:word <= a62[42];
					246:word <= a62[43];
					245:word <= a62[44];
					244:word <= a62[45];
					243:word <= a62[46];
					242:word <= a62[47];
					241:word <= a62[48];
					240:word <= a62[49];
					239:word <= a62[50];
					238:word <= a62[51];
					237:word <= a62[52];
					236:word <= a62[53];
					235:word <= a62[54];
					234:word <= a62[55];
					233:word <= a62[56];
					232:word <= a62[57];
					231:word <= a62[58];
					230:word <= a62[59];
					229:word <= a62[60];
					228:word <= a62[61];
					227:word <= a62[62];
					226:word <= a62[63];
					225:word <= a62[64];
					224:word <= a62[65];
					223:word <= a62[66];
					222:word <= a62[67];
					221:word <= a62[68];
					220:word <= a62[69];
					219:word <= a62[70];
					218:word <= a62[71];
					217:word <= a62[72];
					216:word <= a62[73];
					215:word <= a62[74];
					214:word <= a62[75];
					213:word <= a62[76];
					212:word <= a62[77];
					211:word <= a62[78];
					default:word <= a62[79];
					endcase
				end
				103:begin
				case(x)
					290:word <= a63[0];
					289:word <= a63[1];
					287:word <= a63[2];
					286:word <= a63[3];
					285:word <= a63[4];
					284:word <= a63[5];
					283:word <= a63[6];
					282:word <= a63[7];
					281:word <= a63[8];
					280:word <= a63[9];
					279:word <= a63[10];
					278:word <= a63[11];
					277:word <= a63[12];
					276:word <= a63[13];
					275:word <= a63[14];
					274:word <= a63[15];
					273:word <= a63[16];
					272:word <= a63[17];
					271:word <= a63[18];
					270:word <= a63[19];
					269:word <= a63[20];
					268:word <= a63[21];
					267:word <= a63[22];
					266:word <= a63[23];
					265:word <= a63[24];
					264:word <= a63[25];
					263:word <= a63[26];
					262:word <= a63[27];
					261:word <= a63[28];
					260:word <= a63[29];
					259:word <= a63[30];
					258:word <= a63[31];
					257:word <= a63[32];
					256:word <= a63[33];
					255:word <= a63[34];
					254:word <= a63[35];
					253:word <= a63[36];
					252:word <= a63[37];
					251:word <= a63[38];
					250:word <= a63[39];
					249:word <= a63[40];
					248:word <= a63[41];
					247:word <= a63[42];
					246:word <= a63[43];
					245:word <= a63[44];
					244:word <= a63[45];
					243:word <= a63[46];
					242:word <= a63[47];
					241:word <= a63[48];
					240:word <= a63[49];
					239:word <= a63[50];
					238:word <= a63[51];
					237:word <= a63[52];
					236:word <= a63[53];
					235:word <= a63[54];
					234:word <= a63[55];
					233:word <= a63[56];
					232:word <= a63[57];
					231:word <= a63[58];
					230:word <= a63[59];
					229:word <= a63[60];
					228:word <= a63[61];
					227:word <= a63[62];
					226:word <= a63[63];
					225:word <= a63[64];
					224:word <= a63[65];
					223:word <= a63[66];
					222:word <= a63[67];
					221:word <= a63[68];
					220:word <= a63[69];
					219:word <= a63[70];
					218:word <= a63[71];
					217:word <= a63[72];
					216:word <= a63[74];
					215:word <= a63[73];
					214:word <= a63[75];
					213:word <= a63[76];
					212:word <= a63[77];
					211:word <= a63[78];
					default:word <= a63[79];
					endcase
				end
				104:begin
				case(x)
					290:word <= a64[0];
					289:word <= a64[1];
					287:word <= a64[2];
					286:word <= a64[3];
					285:word <= a64[4];
					284:word <= a64[5];
					283:word <= a64[6];
					282:word <= a64[7];
					281:word <= a64[8];
					280:word <= a64[9];
					279:word <= a64[10];
					278:word <= a64[11];
					277:word <= a64[12];
					276:word <= a64[13];
					275:word <= a64[14];
					274:word <= a64[15];
					273:word <= a64[16];
					272:word <= a64[17];
					271:word <= a64[18];
					270:word <= a64[19];
					269:word <= a64[20];
					268:word <= a64[21];
					267:word <= a64[22];
					266:word <= a64[23];
					265:word <= a64[24];
					264:word <= a64[25];
					263:word <= a64[26];
					262:word <= a64[27];
					261:word <= a64[28];
					260:word <= a64[29];
					259:word <= a64[30];
					258:word <= a64[31];
					257:word <= a64[32];
					256:word <= a64[33];
					255:word <= a64[34];
					254:word <= a64[35];
					253:word <= a64[36];
					252:word <= a64[37];
					251:word <= a64[38];
					250:word <= a64[39];
					249:word <= a64[40];
					248:word <= a64[41];
					247:word <= a64[42];
					246:word <= a64[43];
					245:word <= a64[44];
					244:word <= a64[45];
					243:word <= a64[46];
					242:word <= a64[47];
					241:word <= a64[48];
					240:word <= a64[49];
					239:word <= a64[50];
					238:word <= a64[51];
					237:word <= a64[52];
					236:word <= a64[53];
					235:word <= a64[54];
					234:word <= a64[55];
					233:word <= a64[56];
					232:word <= a64[57];
					231:word <= a64[58];
					230:word <= a64[59];
					229:word <= a64[60];
					228:word <= a64[61];
					227:word <= a64[62];
					226:word <= a64[63];
					225:word <= a64[64];
					224:word <= a64[65];
					223:word <= a64[66];
					222:word <= a64[67];
					221:word <= a64[68];
					220:word <= a64[69];
					219:word <= a64[70];
					218:word <= a64[71];
					217:word <= a64[72];
					216:word <= a64[73];
					215:word <= a64[74];
					214:word <= a64[75];
					213:word <= a64[76];
					212:word <= a64[77];
					211:word <= a64[78];
					default:word <= a64[79];
					endcase
				end
				105:begin
				case(x)
					290:word <= a65[0];
					289:word <= a65[1];
					287:word <= a65[2];
					286:word <= a65[3];
					285:word <= a65[4];
					284:word <= a65[5];
					283:word <= a65[6];
					282:word <= a65[7];
					281:word <= a65[8];
					280:word <= a65[9];
					279:word <= a65[10];
					278:word <= a65[11];
					277:word <= a65[12];
					276:word <= a65[13];
					275:word <= a65[14];
					274:word <= a65[15];
					273:word <= a65[16];
					272:word <= a65[17];
					271:word <= a65[18];
					270:word <= a65[19];
					269:word <= a65[20];
					268:word <= a65[21];
					267:word <= a65[22];
					266:word <= a65[23];
					265:word <= a65[24];
					264:word <= a65[25];
					263:word <= a65[26];
					262:word <= a65[27];
					261:word <= a65[28];
					260:word <= a65[29];
					259:word <= a65[30];
					258:word <= a65[31];
					257:word <= a65[32];
					256:word <= a65[33];
					255:word <= a65[34];
					254:word <= a65[35];
					253:word <= a65[36];
					252:word <= a65[37];
					251:word <= a65[38];
					250:word <= a65[39];
					249:word <= a65[40];
					248:word <= a65[41];
					247:word <= a65[42];
					246:word <= a65[43];
					245:word <= a65[44];
					244:word <= a65[45];
					243:word <= a65[46];
					242:word <= a65[47];
					241:word <= a65[48];
					240:word <= a65[49];
					239:word <= a65[50];
					238:word <= a65[51];
					237:word <= a65[52];
					236:word <= a65[53];
					235:word <= a65[54];
					234:word <= a65[55];
					233:word <= a65[56];
					232:word <= a65[57];
					231:word <= a65[58];
					230:word <= a65[59];
					229:word <= a65[60];
					228:word <= a65[61];
					227:word <= a65[62];
					226:word <= a65[63];
					225:word <= a65[64];
					224:word <= a65[65];
					223:word <= a65[66];
					222:word <= a65[67];
					221:word <= a65[68];
					220:word <= a65[69];
					219:word <= a65[70];
					218:word <= a65[71];
					217:word <= a65[72];
					216:word <= a65[73];
					215:word <= a65[74];
					214:word <= a65[75];
					213:word <= a65[76];
					212:word <= a65[77];
					211:word <= a65[78];
					default:word <= a65[79];
					endcase
				end
				106:begin
				case(x)
					290:word <= a66[0];
					289:word <= a66[1];
					287:word <= a66[2];
					286:word <= a66[3];
					285:word <= a66[4];
					284:word <= a66[5];
					283:word <= a66[6];
					282:word <= a66[7];
					281:word <= a66[8];
					280:word <= a66[9];
					279:word <= a66[10];
					278:word <= a66[11];
					277:word <= a66[12];
					276:word <= a66[13];
					275:word <= a66[14];
					274:word <= a66[15];
					273:word <= a66[16];
					272:word <= a66[17];
					271:word <= a66[18];
					270:word <= a66[19];
					269:word <= a66[20];
					268:word <= a66[21];
					267:word <= a66[22];
					266:word <= a66[23];
					265:word <= a66[24];
					264:word <= a66[25];
					263:word <= a66[26];
					262:word <= a66[27];
					261:word <= a66[28];
					260:word <= a66[29];
					259:word <= a66[30];
					258:word <= a66[31];
					257:word <= a66[32];
					256:word <= a66[33];
					255:word <= a66[34];
					254:word <= a66[35];
					253:word <= a66[36];
					252:word <= a66[37];
					251:word <= a66[38];
					250:word <= a66[39];
					249:word <= a66[40];
					248:word <= a66[41];
					247:word <= a66[42];
					246:word <= a66[43];
					245:word <= a66[44];
					244:word <= a66[45];
					243:word <= a66[46];
					242:word <= a66[47];
					241:word <= a66[48];
					240:word <= a66[49];
					239:word <= a66[50];
					238:word <= a66[51];
					237:word <= a66[52];
					236:word <= a66[53];
					235:word <= a66[54];
					234:word <= a66[55];
					233:word <= a66[56];
					232:word <= a66[57];
					231:word <= a66[58];
					230:word <= a66[59];
					229:word <= a66[60];
					228:word <= a66[61];
					227:word <= a66[62];
					226:word <= a66[63];
					225:word <= a66[64];
					224:word <= a66[65];
					223:word <= a66[66];
					222:word <= a66[67];
					221:word <= a66[68];
					220:word <= a66[69];
					219:word <= a66[70];
					218:word <= a66[71];
					217:word <= a66[72];
					216:word <= a66[73];
					215:word <= a66[74];
					214:word <= a66[75];
					213:word <= a66[76];
					212:word <= a66[77];
					211:word <= a66[78];
					default:word <= a66[79];
					endcase
				end
				107:begin
				case(x)
					290:word <= a67[0];
					289:word <= a67[1];
					287:word <= a67[2];
					286:word <= a67[3];
					285:word <= a67[4];
					284:word <= a67[5];
					283:word <= a67[6];
					282:word <= a67[7];
					281:word <= a67[8];
					280:word <= a67[9];
					279:word <= a67[10];
					278:word <= a67[11];
					277:word <= a67[12];
					276:word <= a67[13];
					275:word <= a67[14];
					274:word <= a67[15];
					273:word <= a67[16];
					272:word <= a67[17];
					271:word <= a67[18];
					270:word <= a67[19];
					269:word <= a67[20];
					268:word <= a67[21];
					267:word <= a67[22];
					266:word <= a67[23];
					265:word <= a67[24];
					264:word <= a67[25];
					263:word <= a67[26];
					262:word <= a67[27];
					261:word <= a67[28];
					260:word <= a67[29];
					259:word <= a67[30];
					258:word <= a67[31];
					257:word <= a67[32];
					256:word <= a67[33];
					255:word <= a67[34];
					254:word <= a67[35];
					253:word <= a67[36];
					252:word <= a67[37];
					251:word <= a67[38];
					250:word <= a67[39];
					249:word <= a67[40];
					248:word <= a67[41];
					247:word <= a67[42];
					246:word <= a67[43];
					245:word <= a67[44];
					244:word <= a67[45];
					243:word <= a67[46];
					242:word <= a67[47];
					241:word <= a67[48];
					240:word <= a67[49];
					239:word <= a67[50];
					238:word <= a67[51];
					237:word <= a67[52];
					236:word <= a67[53];
					235:word <= a67[54];
					234:word <= a67[55];
					233:word <= a67[56];
					232:word <= a67[57];
					231:word <= a67[58];
					230:word <= a67[59];
					229:word <= a67[60];
					228:word <= a67[61];
					227:word <= a67[62];
					226:word <= a67[63];
					225:word <= a67[64];
					224:word <= a67[65];
					223:word <= a67[66];
					222:word <= a67[67];
					221:word <= a67[68];
					220:word <= a67[69];
					219:word <= a67[70];
					218:word <= a67[71];
					217:word <= a67[72];
					216:word <= a67[73];
					215:word <= a67[74];
					214:word <= a67[75];
					213:word <= a67[76];
					212:word <= a67[77];
					211:word <= a67[78];
					default:word <= a67[79];
					endcase
				end
				108:begin
				case(x)
					290:word <= a68[0];
					289:word <= a68[1];
					287:word <= a68[2];
					286:word <= a68[3];
					285:word <= a68[4];
					284:word <= a68[5];
					283:word <= a68[6];
					282:word <= a68[7];
					281:word <= a68[8];
					280:word <= a68[9];
					279:word <= a68[10];
					278:word <= a68[11];
					277:word <= a68[12];
					276:word <= a68[13];
					275:word <= a68[14];
					274:word <= a68[15];
					273:word <= a68[16];
					272:word <= a68[17];
					271:word <= a68[18];
					270:word <= a68[19];
					269:word <= a68[20];
					268:word <= a68[21];
					267:word <= a68[22];
					266:word <= a68[23];
					265:word <= a68[24];
					264:word <= a68[25];
					263:word <= a68[26];
					262:word <= a68[27];
					261:word <= a68[28];
					260:word <= a68[29];
					259:word <= a68[30];
					258:word <= a68[31];
					257:word <= a68[32];
					256:word <= a68[33];
					255:word <= a68[34];
					254:word <= a68[35];
					253:word <= a68[36];
					252:word <= a68[37];
					251:word <= a68[38];
					250:word <= a68[39];
					249:word <= a68[40];
					248:word <= a68[41];
					247:word <= a68[42];
					246:word <= a68[43];
					245:word <= a68[44];
					244:word <= a68[45];
					243:word <= a68[46];
					242:word <= a68[47];
					241:word <= a68[48];
					240:word <= a68[49];
					239:word <= a68[50];
					238:word <= a68[51];
					237:word <= a68[52];
					236:word <= a68[53];
					235:word <= a68[54];
					234:word <= a68[55];
					233:word <= a68[56];
					232:word <= a68[57];
					231:word <= a68[58];
					230:word <= a68[59];
					229:word <= a68[60];
					228:word <= a68[61];
					227:word <= a68[62];
					226:word <= a68[63];
					225:word <= a68[64];
					224:word <= a68[65];
					223:word <= a68[66];
					222:word <= a68[67];
					221:word <= a68[68];
					220:word <= a68[69];
					219:word <= a68[70];
					218:word <= a68[71];
					217:word <= a68[72];
					216:word <= a68[73];
					215:word <= a68[74];
					214:word <= a68[75];
					213:word <= a68[76];
					212:word <= a68[77];
					211:word <= a68[78];
					default:word <= a68[79];
					endcase
				end
				109:begin
				case(x)
					290:word <= a69[0];
					289:word <= a69[1];
					287:word <= a69[2];
					286:word <= a69[3];
					285:word <= a69[4];
					284:word <= a69[5];
					283:word <= a69[6];
					282:word <= a69[7];
					281:word <= a69[8];
					280:word <= a69[9];
					279:word <= a69[10];
					278:word <= a69[11];
					277:word <= a69[12];
					276:word <= a69[13];
					275:word <= a69[14];
					274:word <= a69[15];
					273:word <= a69[16];
					272:word <= a69[17];
					271:word <= a69[18];
					270:word <= a69[19];
					269:word <= a69[20];
					268:word <= a69[21];
					267:word <= a69[22];
					266:word <= a69[23];
					265:word <= a69[24];
					264:word <= a69[25];
					263:word <= a69[26];
					262:word <= a69[27];
					261:word <= a69[28];
					260:word <= a69[29];
					259:word <= a69[30];
					258:word <= a69[31];
					257:word <= a69[32];
					256:word <= a69[33];
					255:word <= a69[34];
					254:word <= a69[35];
					253:word <= a69[36];
					252:word <= a69[37];
					251:word <= a69[38];
					250:word <= a69[39];
					249:word <= a69[40];
					248:word <= a69[41];
					247:word <= a69[42];
					246:word <= a69[43];
					245:word <= a69[44];
					244:word <= a69[45];
					243:word <= a69[46];
					242:word <= a69[47];
					241:word <= a69[48];
					240:word <= a69[49];
					239:word <= a69[50];
					238:word <= a69[51];
					237:word <= a69[52];
					236:word <= a69[53];
					235:word <= a69[54];
					234:word <= a69[55];
					233:word <= a69[56];
					232:word <= a69[57];
					231:word <= a69[58];
					230:word <= a69[59];
					229:word <= a69[60];
					228:word <= a69[61];
					227:word <= a69[62];
					226:word <= a69[63];
					225:word <= a69[64];
					224:word <= a69[65];
					223:word <= a69[66];
					222:word <= a69[67];
					221:word <= a69[68];
					220:word <= a69[69];
					219:word <= a69[70];
					218:word <= a69[71];
					217:word <= a69[72];
					216:word <= a69[73];
					215:word <= a69[74];
					214:word <= a69[75];
					213:word <= a69[76];
					212:word <= a69[77];
					211:word <= a69[78];
					default:word <= a69[79];
					endcase
				end
				110:begin
				case(x)
					290:word <= a70[0];
					289:word <= a70[1];
					287:word <= a70[2];
					286:word <= a70[3];
					285:word <= a70[4];
					284:word <= a70[5];
					283:word <= a70[6];
					282:word <= a70[7];
					281:word <= a70[8];
					280:word <= a70[9];
					279:word <= a70[10];
					278:word <= a70[11];
					277:word <= a70[12];
					276:word <= a70[13];
					275:word <= a70[14];
					274:word <= a70[15];
					273:word <= a70[16];
					272:word <= a70[17];
					271:word <= a70[18];
					270:word <= a70[19];
					269:word <= a70[20];
					268:word <= a70[21];
					267:word <= a70[22];
					266:word <= a70[23];
					265:word <= a70[24];
					264:word <= a70[25];
					263:word <= a70[26];
					262:word <= a70[27];
					261:word <= a70[28];
					260:word <= a70[29];
					259:word <= a70[30];
					258:word <= a70[31];
					257:word <= a70[32];
					256:word <= a70[33];
					255:word <= a70[34];
					254:word <= a70[35];
					253:word <= a70[36];
					252:word <= a70[37];
					251:word <= a70[38];
					250:word <= a70[39];
					249:word <= a70[40];
					248:word <= a70[41];
					247:word <= a70[42];
					246:word <= a70[43];
					245:word <= a70[44];
					244:word <= a70[45];
					243:word <= a70[46];
					242:word <= a70[47];
					241:word <= a70[48];
					240:word <= a70[49];
					239:word <= a70[50];
					238:word <= a70[51];
					237:word <= a70[52];
					236:word <= a70[53];
					235:word <= a70[54];
					234:word <= a70[55];
					233:word <= a70[56];
					232:word <= a70[57];
					231:word <= a70[58];
					230:word <= a70[59];
					229:word <= a70[60];
					228:word <= a70[61];
					227:word <= a70[62];
					226:word <= a70[63];
					225:word <= a70[64];
					224:word <= a70[65];
					223:word <= a70[66];
					222:word <= a70[67];
					221:word <= a70[68];
					220:word <= a70[69];
					219:word <= a70[70];
					218:word <= a70[71];
					217:word <= a70[72];
					216:word <= a70[73];
					215:word <= a70[74];
					214:word <= a70[75];
					213:word <= a70[76];
					212:word <= a70[77];
					211:word <= a70[78];
					default:word <= a70[79];
					endcase
				end
				111:begin
				case(x)
					290:word <= a71[0];
					289:word <= a71[1];
					287:word <= a71[2];
					286:word <= a71[3];
					285:word <= a71[4];
					284:word <= a71[5];
					283:word <= a71[6];
					282:word <= a71[7];
					281:word <= a71[8];
					280:word <= a71[9];
					279:word <= a71[10];
					278:word <= a71[11];
					277:word <= a71[12];
					276:word <= a71[13];
					275:word <= a71[14];
					274:word <= a71[15];
					273:word <= a71[16];
					272:word <= a71[17];
					271:word <= a71[18];
					270:word <= a71[19];
					269:word <= a71[20];
					268:word <= a71[21];
					267:word <= a71[22];
					266:word <= a71[23];
					265:word <= a71[24];
					264:word <= a71[25];
					263:word <= a71[26];
					262:word <= a71[27];
					261:word <= a71[28];
					260:word <= a71[29];
					259:word <= a71[30];
					258:word <= a71[31];
					257:word <= a71[32];
					256:word <= a71[33];
					255:word <= a71[34];
					254:word <= a71[35];
					253:word <= a71[36];
					252:word <= a71[37];
					251:word <= a71[38];
					250:word <= a71[39];
					249:word <= a71[40];
					248:word <= a71[41];
					247:word <= a71[42];
					246:word <= a71[43];
					245:word <= a71[44];
					244:word <= a71[45];
					243:word <= a71[46];
					242:word <= a71[47];
					241:word <= a71[48];
					240:word <= a71[49];
					239:word <= a71[50];
					238:word <= a71[51];
					237:word <= a71[52];
					236:word <= a71[53];
					235:word <= a71[54];
					234:word <= a71[55];
					233:word <= a71[56];
					232:word <= a71[57];
					231:word <= a71[58];
					230:word <= a71[59];
					229:word <= a71[60];
					228:word <= a71[61];
					227:word <= a71[62];
					226:word <= a71[63];
					225:word <= a71[64];
					224:word <= a71[65];
					223:word <= a71[66];
					222:word <= a71[67];
					221:word <= a71[68];
					220:word <= a71[69];
					219:word <= a71[70];
					218:word <= a71[71];
					217:word <= a71[72];
					216:word <= a71[73];
					215:word <= a71[74];
					214:word <= a71[75];
					213:word <= a71[76];
					212:word <= a71[77];
					211:word <= a71[78];
					default:word <= a71[79];
					endcase
				end
				112:begin
				case(x)
					290:word <= a72[0];
					289:word <= a72[1];
					287:word <= a72[2];
					286:word <= a72[3];
					285:word <= a72[4];
					284:word <= a72[5];
					283:word <= a72[6];
					282:word <= a72[7];
					281:word <= a72[8];
					280:word <= a72[9];
					279:word <= a72[10];
					278:word <= a72[11];
					277:word <= a72[12];
					276:word <= a72[13];
					275:word <= a72[14];
					274:word <= a72[15];
					273:word <= a72[16];
					272:word <= a72[17];
					271:word <= a72[18];
					270:word <= a72[19];
					269:word <= a72[20];
					268:word <= a72[21];
					267:word <= a72[22];
					266:word <= a72[23];
					265:word <= a72[24];
					264:word <= a72[25];
					263:word <= a72[26];
					262:word <= a72[27];
					261:word <= a72[28];
					260:word <= a72[29];
					259:word <= a72[30];
					258:word <= a72[31];
					257:word <= a72[32];
					256:word <= a72[33];
					255:word <= a72[34];
					254:word <= a72[35];
					253:word <= a72[36];
					252:word <= a72[37];
					251:word <= a72[38];
					250:word <= a72[39];
					249:word <= a72[40];
					248:word <= a72[41];
					247:word <= a72[42];
					246:word <= a72[43];
					245:word <= a72[44];
					244:word <= a72[45];
					243:word <= a72[46];
					242:word <= a72[47];
					241:word <= a72[48];
					240:word <= a72[49];
					239:word <= a72[50];
					238:word <= a72[51];
					237:word <= a72[52];
					236:word <= a72[53];
					235:word <= a72[54];
					234:word <= a72[55];
					233:word <= a72[56];
					232:word <= a72[57];
					231:word <= a72[58];
					230:word <= a72[59];
					229:word <= a72[60];
					228:word <= a72[61];
					227:word <= a72[62];
					226:word <= a72[63];
					225:word <= a72[64];
					224:word <= a72[65];
					223:word <= a72[66];
					222:word <= a72[67];
					221:word <= a72[68];
					220:word <= a72[69];
					219:word <= a72[70];
					218:word <= a72[71];
					217:word <= a72[72];
					216:word <= a72[73];
					215:word <= a72[74];
					214:word <= a72[75];
					213:word <= a72[76];
					212:word <= a72[77];
					211:word <= a72[78];
					default:word <= a72[79];
					endcase
				end
				113:begin
				case(x)
					290:word <= a73[0];
					289:word <= a73[1];
					287:word <= a73[2];
					286:word <= a73[3];
					285:word <= a73[4];
					284:word <= a73[5];
					283:word <= a73[6];
					282:word <= a73[7];
					281:word <= a73[8];
					280:word <= a73[9];
					279:word <= a73[10];
					278:word <= a73[11];
					277:word <= a73[12];
					276:word <= a73[13];
					275:word <= a73[14];
					274:word <= a73[15];
					273:word <= a73[16];
					272:word <= a73[17];
					271:word <= a73[18];
					270:word <= a73[19];
					269:word <= a73[20];
					268:word <= a73[21];
					267:word <= a73[22];
					266:word <= a73[23];
					265:word <= a73[24];
					264:word <= a73[25];
					263:word <= a73[26];
					262:word <= a73[27];
					261:word <= a73[28];
					260:word <= a73[29];
					259:word <= a73[30];
					258:word <= a73[31];
					257:word <= a73[32];
					256:word <= a73[33];
					255:word <= a73[34];
					254:word <= a73[35];
					253:word <= a73[36];
					252:word <= a73[37];
					251:word <= a73[38];
					250:word <= a73[39];
					249:word <= a73[40];
					248:word <= a73[41];
					247:word <= a73[42];
					246:word <= a73[43];
					245:word <= a73[44];
					244:word <= a73[45];
					243:word <= a73[46];
					242:word <= a73[47];
					241:word <= a73[48];
					240:word <= a73[49];
					239:word <= a73[50];
					238:word <= a73[51];
					237:word <= a73[52];
					236:word <= a73[53];
					235:word <= a73[54];
					234:word <= a73[55];
					233:word <= a73[56];
					232:word <= a73[57];
					231:word <= a73[58];
					230:word <= a73[59];
					229:word <= a73[60];
					228:word <= a73[61];
					227:word <= a73[62];
					226:word <= a73[63];
					225:word <= a73[64];
					224:word <= a73[65];
					223:word <= a73[66];
					222:word <= a73[67];
					221:word <= a73[68];
					220:word <= a73[69];
					219:word <= a73[70];
					218:word <= a73[71];
					217:word <= a73[72];
					216:word <= a73[73];
					215:word <= a73[74];
					214:word <= a73[75];
					213:word <= a73[76];
					212:word <= a73[77];
					211:word <= a73[78];
					default:word <= a73[79];
					endcase
				end
				114:begin
				case(x)
					290:word <= a74[0];
					289:word <= a74[1];
					287:word <= a74[2];
					286:word <= a74[3];
					285:word <= a74[4];
					284:word <= a74[5];
					283:word <= a74[6];
					282:word <= a74[7];
					281:word <= a74[8];
					280:word <= a74[9];
					279:word <= a74[10];
					278:word <= a74[11];
					277:word <= a74[12];
					276:word <= a74[13];
					275:word <= a74[14];
					274:word <= a74[15];
					273:word <= a74[16];
					272:word <= a74[17];
					271:word <= a74[18];
					270:word <= a74[19];
					269:word <= a74[20];
					268:word <= a74[21];
					267:word <= a74[22];
					266:word <= a74[23];
					265:word <= a74[24];
					264:word <= a74[25];
					263:word <= a74[26];
					262:word <= a74[27];
					261:word <= a74[28];
					260:word <= a74[29];
					259:word <= a74[30];
					258:word <= a74[31];
					257:word <= a74[32];
					256:word <= a74[33];
					255:word <= a74[34];
					254:word <= a74[35];
					253:word <= a74[36];
					252:word <= a74[37];
					251:word <= a74[38];
					250:word <= a74[39];
					249:word <= a74[40];
					248:word <= a74[41];
					247:word <= a74[42];
					246:word <= a74[43];
					245:word <= a74[44];
					244:word <= a74[45];
					243:word <= a74[46];
					242:word <= a74[47];
					241:word <= a74[48];
					240:word <= a74[49];
					239:word <= a74[50];
					238:word <= a74[51];
					237:word <= a74[52];
					236:word <= a74[53];
					235:word <= a74[54];
					234:word <= a74[55];
					233:word <= a74[56];
					232:word <= a74[57];
					231:word <= a74[58];
					230:word <= a74[59];
					229:word <= a74[60];
					228:word <= a74[61];
					227:word <= a74[62];
					226:word <= a74[63];
					225:word <= a74[64];
					224:word <= a74[65];
					223:word <= a74[66];
					222:word <= a74[67];
					221:word <= a74[68];
					220:word <= a74[69];
					219:word <= a74[70];
					218:word <= a74[71];
					217:word <= a74[72];
					216:word <= a74[73];
					215:word <= a74[74];
					214:word <= a74[75];
					213:word <= a74[76];
					212:word <= a74[77];
					211:word <= a74[78];
					default:word <= a74[79];
					endcase
				end
				115:begin
				case(x)
					290:word <= a75[0];
					289:word <= a75[1];
					287:word <= a75[2];
					286:word <= a75[3];
					285:word <= a75[4];
					284:word <= a75[5];
					283:word <= a75[6];
					282:word <= a75[7];
					281:word <= a75[8];
					280:word <= a75[9];
					279:word <= a75[10];
					278:word <= a75[11];
					277:word <= a75[12];
					276:word <= a75[13];
					275:word <= a75[14];
					274:word <= a75[15];
					273:word <= a75[16];
					272:word <= a75[17];
					271:word <= a75[18];
					270:word <= a75[19];
					269:word <= a75[20];
					268:word <= a75[21];
					267:word <= a75[22];
					266:word <= a75[23];
					265:word <= a75[24];
					264:word <= a75[25];
					263:word <= a75[26];
					262:word <= a75[27];
					261:word <= a75[28];
					260:word <= a75[29];
					259:word <= a75[30];
					258:word <= a75[31];
					257:word <= a75[32];
					256:word <= a75[33];
					255:word <= a75[34];
					254:word <= a75[35];
					253:word <= a75[36];
					252:word <= a75[37];
					251:word <= a75[38];
					250:word <= a75[39];
					249:word <= a75[40];
					248:word <= a75[41];
					247:word <= a75[42];
					246:word <= a75[43];
					245:word <= a75[44];
					244:word <= a75[45];
					243:word <= a75[46];
					242:word <= a75[47];
					241:word <= a75[48];
					240:word <= a75[49];
					239:word <= a75[50];
					238:word <= a75[51];
					237:word <= a75[52];
					236:word <= a75[53];
					235:word <= a75[54];
					234:word <= a75[55];
					233:word <= a75[56];
					232:word <= a75[57];
					231:word <= a75[58];
					230:word <= a75[59];
					229:word <= a75[60];
					228:word <= a75[61];
					227:word <= a75[62];
					226:word <= a75[63];
					225:word <= a75[64];
					224:word <= a75[65];
					223:word <= a75[66];
					222:word <= a75[67];
					221:word <= a75[68];
					220:word <= a75[69];
					219:word <= a75[70];
					218:word <= a75[71];
					217:word <= a75[72];
					216:word <= a75[73];
					215:word <= a75[74];
					214:word <= a75[75];
					213:word <= a75[76];
					212:word <= a75[77];
					211:word <= a75[78];
					default:word <= a75[79];
					endcase
				end
				116:begin
				case(x)
					290:word <= a76[0];
					289:word <= a76[1];
					287:word <= a76[2];
					286:word <= a76[3];
					285:word <= a76[4];
					284:word <= a76[5];
					283:word <= a76[6];
					282:word <= a76[7];
					281:word <= a76[8];
					280:word <= a76[9];
					279:word <= a76[10];
					278:word <= a76[11];
					277:word <= a76[12];
					276:word <= a76[13];
					275:word <= a76[14];
					274:word <= a76[15];
					273:word <= a76[16];
					272:word <= a76[17];
					271:word <= a76[18];
					270:word <= a76[19];
					269:word <= a76[20];
					268:word <= a76[21];
					267:word <= a76[22];
					266:word <= a76[23];
					265:word <= a76[24];
					264:word <= a76[25];
					263:word <= a76[26];
					262:word <= a76[27];
					261:word <= a76[28];
					260:word <= a76[29];
					259:word <= a76[30];
					258:word <= a76[31];
					257:word <= a76[32];
					256:word <= a76[33];
					255:word <= a76[34];
					254:word <= a76[35];
					253:word <= a76[36];
					252:word <= a76[37];
					251:word <= a76[38];
					250:word <= a76[39];
					249:word <= a76[40];
					248:word <= a76[41];
					247:word <= a76[42];
					246:word <= a76[43];
					245:word <= a76[44];
					244:word <= a76[45];
					243:word <= a76[46];
					242:word <= a76[47];
					241:word <= a76[48];
					240:word <= a76[49];
					239:word <= a76[50];
					238:word <= a76[51];
					237:word <= a76[52];
					236:word <= a76[53];
					235:word <= a76[54];
					234:word <= a76[55];
					233:word <= a76[56];
					232:word <= a76[57];
					231:word <= a76[58];
					230:word <= a76[59];
					229:word <= a76[60];
					228:word <= a76[61];
					227:word <= a76[62];
					226:word <= a76[63];
					225:word <= a76[64];
					224:word <= a76[65];
					223:word <= a76[66];
					222:word <= a76[67];
					221:word <= a76[68];
					220:word <= a76[69];
					219:word <= a76[70];
					218:word <= a76[71];
					217:word <= a76[72];
					216:word <= a76[73];
					215:word <= a76[74];
					214:word <= a76[75];
					213:word <= a76[76];
					212:word <= a76[77];
					211:word <= a76[78];
					default:word <= a76[79];
					endcase
				end
				117:begin
				case(x)
					290:word <= a77[0];
					289:word <= a77[1];
					287:word <= a77[2];
					286:word <= a77[3];
					285:word <= a77[4];
					284:word <= a77[5];
					283:word <= a77[6];
					282:word <= a77[7];
					281:word <= a77[8];
					280:word <= a77[9];
					279:word <= a77[10];
					278:word <= a77[11];
					277:word <= a77[12];
					276:word <= a77[13];
					275:word <= a77[14];
					274:word <= a77[15];
					273:word <= a77[16];
					272:word <= a77[17];
					271:word <= a77[18];
					270:word <= a77[19];
					269:word <= a77[20];
					268:word <= a77[21];
					267:word <= a77[22];
					266:word <= a77[23];
					265:word <= a77[24];
					264:word <= a77[25];
					263:word <= a77[26];
					262:word <= a77[27];
					261:word <= a77[28];
					260:word <= a77[29];
					259:word <= a77[30];
					258:word <= a77[31];
					257:word <= a77[32];
					256:word <= a77[33];
					255:word <= a77[34];
					254:word <= a77[35];
					253:word <= a77[36];
					252:word <= a77[37];
					251:word <= a77[38];
					250:word <= a77[39];
					249:word <= a77[40];
					248:word <= a77[41];
					247:word <= a77[42];
					246:word <= a77[43];
					245:word <= a77[44];
					244:word <= a77[45];
					243:word <= a77[46];
					242:word <= a77[47];
					241:word <= a77[48];
					240:word <= a77[49];
					239:word <= a77[50];
					238:word <= a77[51];
					237:word <= a77[52];
					236:word <= a77[53];
					235:word <= a77[54];
					234:word <= a77[55];
					233:word <= a77[56];
					232:word <= a77[57];
					231:word <= a77[58];
					230:word <= a77[59];
					229:word <= a77[60];
					228:word <= a77[61];
					227:word <= a77[62];
					226:word <= a77[63];
					225:word <= a77[64];
					224:word <= a77[65];
					223:word <= a77[66];
					222:word <= a77[67];
					221:word <= a77[68];
					220:word <= a77[69];
					219:word <= a77[70];
					218:word <= a77[71];
					217:word <= a77[72];
					216:word <= a77[73];
					215:word <= a77[74];
					214:word <= a77[75];
					213:word <= a77[76];
					212:word <= a77[77];
					211:word <= a77[78];
					default:word <= a77[79];
					endcase
				end
				118:begin
				case(x)
					290:word <= a78[0];
					289:word <= a78[1];
					287:word <= a78[2];
					286:word <= a78[3];
					285:word <= a78[4];
					284:word <= a78[5];
					283:word <= a78[6];
					282:word <= a78[7];
					281:word <= a78[8];
					280:word <= a78[9];
					279:word <= a78[10];
					278:word <= a78[11];
					277:word <= a78[12];
					276:word <= a78[13];
					275:word <= a78[14];
					274:word <= a78[15];
					273:word <= a78[16];
					272:word <= a78[17];
					271:word <= a78[18];
					270:word <= a78[19];
					269:word <= a78[20];
					268:word <= a78[21];
					267:word <= a78[22];
					266:word <= a78[23];
					265:word <= a78[24];
					264:word <= a78[25];
					263:word <= a78[26];
					262:word <= a78[27];
					261:word <= a78[28];
					260:word <= a78[29];
					259:word <= a78[30];
					258:word <= a78[31];
					257:word <= a78[32];
					256:word <= a78[33];
					255:word <= a78[34];
					254:word <= a78[35];
					253:word <= a78[36];
					252:word <= a78[37];
					251:word <= a78[38];
					250:word <= a78[39];
					249:word <= a78[40];
					248:word <= a78[41];
					247:word <= a78[42];
					246:word <= a78[43];
					245:word <= a78[44];
					244:word <= a78[45];
					243:word <= a78[46];
					242:word <= a78[47];
					241:word <= a78[48];
					240:word <= a78[49];
					239:word <= a78[50];
					238:word <= a78[51];
					237:word <= a78[52];
					236:word <= a78[53];
					235:word <= a78[54];
					234:word <= a78[55];
					233:word <= a78[56];
					232:word <= a78[57];
					231:word <= a78[58];
					230:word <= a78[59];
					229:word <= a78[60];
					228:word <= a78[61];
					227:word <= a78[62];
					226:word <= a78[63];
					225:word <= a78[64];
					224:word <= a78[65];
					223:word <= a78[66];
					222:word <= a78[67];
					221:word <= a78[68];
					220:word <= a78[69];
					219:word <= a78[70];
					218:word <= a78[71];
					217:word <= a78[72];
					216:word <= a78[73];
					215:word <= a78[74];
					214:word <= a78[75];
					213:word <= a78[76];
					212:word <= a78[77];
					211:word <= a78[78];
					default:word <= a78[79];
					endcase
				end
				119:begin
				case(x)
					290:word <= a79[0];
					289:word <= a79[1];
					287:word <= a79[2];
					286:word <= a79[3];
					285:word <= a79[4];
					284:word <= a79[5];
					283:word <= a79[6];
					282:word <= a79[7];
					281:word <= a79[8];
					280:word <= a79[9];
					279:word <= a79[10];
					278:word <= a79[11];
					277:word <= a79[12];
					276:word <= a79[13];
					275:word <= a79[14];
					274:word <= a79[15];
					273:word <= a79[16];
					272:word <= a79[17];
					271:word <= a79[18];
					270:word <= a79[19];
					269:word <= a79[20];
					268:word <= a79[21];
					267:word <= a79[22];
					266:word <= a79[23];
					265:word <= a79[24];
					264:word <= a79[25];
					263:word <= a79[26];
					262:word <= a79[27];
					261:word <= a79[28];
					260:word <= a79[29];
					259:word <= a79[30];
					258:word <= a79[31];
					257:word <= a79[32];
					256:word <= a79[33];
					255:word <= a79[34];
					254:word <= a79[35];
					253:word <= a79[36];
					252:word <= a79[37];
					251:word <= a79[38];
					250:word <= a79[39];
					249:word <= a79[40];
					248:word <= a79[41];
					247:word <= a79[42];
					246:word <= a79[43];
					245:word <= a79[44];
					244:word <= a79[45];
					243:word <= a79[46];
					242:word <= a79[47];
					241:word <= a79[48];
					240:word <= a79[49];
					239:word <= a79[50];
					238:word <= a79[51];
					237:word <= a79[52];
					236:word <= a79[53];
					235:word <= a79[54];
					234:word <= a79[55];
					233:word <= a79[56];
					232:word <= a79[57];
					231:word <= a79[58];
					230:word <= a79[59];
					229:word <= a79[60];
					228:word <= a79[61];
					227:word <= a79[62];
					226:word <= a79[63];
					225:word <= a79[64];
					224:word <= a79[65];
					223:word <= a79[66];
					222:word <= a79[67];
					221:word <= a79[68];
					220:word <= a79[69];
					219:word <= a79[70];
					218:word <= a79[71];
					217:word <= a79[72];
					216:word <= a79[73];
					215:word <= a79[74];
					214:word <= a79[75];
					213:word <= a79[76];
					212:word <= a79[77];
					211:word <= a79[78];
					default:word <= a79[79];
					endcase
				end
				120:begin
				case(x)
					290:word <= a80[0];
					289:word <= a80[1];
					287:word <= a80[2];
					286:word <= a80[3];
					285:word <= a80[4];
					284:word <= a80[5];
					283:word <= a80[6];
					282:word <= a80[7];
					281:word <= a80[8];
					280:word <= a80[9];
					279:word <= a80[10];
					278:word <= a80[11];
					277:word <= a80[12];
					276:word <= a80[13];
					275:word <= a80[14];
					274:word <= a80[15];
					273:word <= a80[16];
					272:word <= a80[17];
					271:word <= a80[18];
					270:word <= a80[19];
					269:word <= a80[20];
					268:word <= a80[21];
					267:word <= a80[22];
					266:word <= a80[23];
					265:word <= a80[24];
					264:word <= a80[25];
					263:word <= a80[26];
					262:word <= a80[27];
					261:word <= a80[28];
					260:word <= a80[29];
					259:word <= a80[30];
					258:word <= a80[31];
					257:word <= a80[32];
					256:word <= a80[33];
					255:word <= a80[34];
					254:word <= a80[35];
					253:word <= a80[36];
					252:word <= a80[37];
					251:word <= a80[38];
					250:word <= a80[39];
					249:word <= a80[40];
					248:word <= a80[41];
					247:word <= a80[42];
					246:word <= a80[43];
					245:word <= a80[44];
					244:word <= a80[45];
					243:word <= a80[46];
					242:word <= a80[47];
					241:word <= a80[48];
					240:word <= a80[49];
					239:word <= a80[50];
					238:word <= a80[51];
					237:word <= a80[52];
					236:word <= a80[53];
					235:word <= a80[54];
					234:word <= a80[55];
					233:word <= a80[56];
					232:word <= a80[57];
					231:word <= a80[58];
					230:word <= a80[59];
					229:word <= a80[60];
					228:word <= a80[61];
					227:word <= a80[62];
					226:word <= a80[63];
					225:word <= a80[64];
					224:word <= a80[65];
					223:word <= a80[66];
					222:word <= a80[67];
					221:word <= a80[68];
					220:word <= a80[69];
					219:word <= a80[70];
					218:word <= a80[71];
					217:word <= a80[72];
					216:word <= a80[73];
					215:word <= a80[74];
					214:word <= a80[75];
					213:word <= a80[76];
					212:word <= a80[77];
					211:word <= a80[78];
					default:word <= a80[79];
					endcase
				end
				121:begin
				case(x)
					290:word <= a81[0];
					289:word <= a81[1];
					287:word <= a81[2];
					286:word <= a81[3];
					285:word <= a81[4];
					284:word <= a81[5];
					283:word <= a81[6];
					282:word <= a81[7];
					281:word <= a81[8];
					280:word <= a81[9];
					279:word <= a81[10];
					278:word <= a81[11];
					277:word <= a81[12];
					276:word <= a81[13];
					275:word <= a81[14];
					274:word <= a81[15];
					273:word <= a81[16];
					272:word <= a81[17];
					271:word <= a81[18];
					270:word <= a81[19];
					269:word <= a81[20];
					268:word <= a81[21];
					267:word <= a81[22];
					266:word <= a81[23];
					265:word <= a81[24];
					264:word <= a81[25];
					263:word <= a81[26];
					262:word <= a81[27];
					261:word <= a81[28];
					260:word <= a81[29];
					259:word <= a81[30];
					258:word <= a81[31];
					257:word <= a81[32];
					256:word <= a81[33];
					255:word <= a81[34];
					254:word <= a81[35];
					253:word <= a81[36];
					252:word <= a81[37];
					251:word <= a81[38];
					250:word <= a81[39];
					249:word <= a81[40];
					248:word <= a81[41];
					247:word <= a81[42];
					246:word <= a81[43];
					245:word <= a81[44];
					244:word <= a81[45];
					243:word <= a81[46];
					242:word <= a81[47];
					241:word <= a81[48];
					240:word <= a81[49];
					239:word <= a81[50];
					238:word <= a81[51];
					237:word <= a81[52];
					236:word <= a81[53];
					235:word <= a81[54];
					234:word <= a81[55];
					233:word <= a81[56];
					232:word <= a81[57];
					231:word <= a81[58];
					230:word <= a81[59];
					229:word <= a81[60];
					228:word <= a81[61];
					227:word <= a81[62];
					226:word <= a81[63];
					225:word <= a81[64];
					224:word <= a81[65];
					223:word <= a81[66];
					222:word <= a81[67];
					221:word <= a81[68];
					220:word <= a81[69];
					219:word <= a81[70];
					218:word <= a81[71];
					217:word <= a81[72];
					216:word <= a81[73];
					215:word <= a81[74];
					214:word <= a81[75];
					213:word <= a81[76];
					212:word <= a81[77];
					211:word <= a81[78];
					default:word <= a81[79];
					endcase
				end
				122:begin
				case(x)
					290:word <= a82[0];
					289:word <= a82[1];
					287:word <= a82[2];
					286:word <= a82[3];
					285:word <= a82[4];
					284:word <= a82[5];
					283:word <= a82[6];
					282:word <= a82[7];
					281:word <= a82[8];
					280:word <= a82[9];
					279:word <= a82[10];
					278:word <= a82[11];
					277:word <= a82[12];
					276:word <= a82[13];
					275:word <= a82[14];
					274:word <= a82[15];
					273:word <= a82[16];
					272:word <= a82[17];
					271:word <= a82[18];
					270:word <= a82[19];
					269:word <= a82[20];
					268:word <= a82[21];
					267:word <= a82[22];
					266:word <= a82[23];
					265:word <= a82[24];
					264:word <= a82[25];
					263:word <= a82[26];
					262:word <= a82[27];
					261:word <= a82[28];
					260:word <= a82[29];
					259:word <= a82[30];
					258:word <= a82[31];
					257:word <= a82[32];
					256:word <= a82[33];
					255:word <= a82[34];
					254:word <= a82[35];
					253:word <= a82[36];
					252:word <= a82[37];
					251:word <= a82[38];
					250:word <= a82[39];
					249:word <= a82[40];
					248:word <= a82[41];
					247:word <= a82[42];
					246:word <= a82[43];
					245:word <= a82[44];
					244:word <= a82[45];
					243:word <= a82[46];
					242:word <= a82[47];
					241:word <= a82[48];
					240:word <= a82[49];
					239:word <= a82[50];
					238:word <= a82[51];
					237:word <= a82[52];
					236:word <= a82[53];
					235:word <= a82[54];
					234:word <= a82[55];
					233:word <= a82[56];
					232:word <= a82[57];
					231:word <= a82[58];
					230:word <= a82[59];
					229:word <= a82[60];
					228:word <= a82[61];
					227:word <= a82[62];
					226:word <= a82[63];
					225:word <= a82[64];
					224:word <= a82[65];
					223:word <= a82[66];
					222:word <= a82[67];
					221:word <= a82[68];
					220:word <= a82[69];
					219:word <= a82[70];
					218:word <= a82[71];
					217:word <= a82[72];
					216:word <= a82[73];
					215:word <= a82[74];
					214:word <= a82[75];
					213:word <= a82[76];
					212:word <= a82[77];
					211:word <= a82[78];
					default:word <= a82[79];
					endcase
				end
				123:begin
				case(x)
					290:word <= a83[0];
					289:word <= a83[1];
					287:word <= a83[2];
					286:word <= a83[3];
					285:word <= a83[4];
					284:word <= a83[5];
					283:word <= a83[6];
					282:word <= a83[7];
					281:word <= a83[8];
					280:word <= a83[9];
					279:word <= a83[10];
					278:word <= a83[11];
					277:word <= a83[12];
					276:word <= a83[13];
					275:word <= a83[14];
					274:word <= a83[15];
					273:word <= a83[16];
					272:word <= a83[17];
					271:word <= a83[18];
					270:word <= a83[19];
					269:word <= a83[20];
					268:word <= a83[21];
					267:word <= a83[22];
					266:word <= a83[23];
					265:word <= a83[24];
					264:word <= a83[25];
					263:word <= a83[26];
					262:word <= a83[27];
					261:word <= a83[28];
					260:word <= a83[29];
					259:word <= a83[30];
					258:word <= a83[31];
					257:word <= a83[32];
					256:word <= a83[33];
					255:word <= a83[34];
					254:word <= a83[35];
					253:word <= a83[36];
					252:word <= a83[37];
					251:word <= a83[38];
					250:word <= a83[39];
					249:word <= a83[40];
					248:word <= a83[41];
					247:word <= a83[42];
					246:word <= a83[43];
					245:word <= a83[44];
					244:word <= a83[45];
					243:word <= a83[46];
					242:word <= a83[47];
					241:word <= a83[48];
					240:word <= a83[49];
					239:word <= a83[50];
					238:word <= a83[51];
					237:word <= a83[52];
					236:word <= a83[53];
					235:word <= a83[54];
					234:word <= a83[55];
					233:word <= a83[56];
					232:word <= a83[57];
					231:word <= a83[58];
					230:word <= a83[59];
					229:word <= a83[60];
					228:word <= a83[61];
					227:word <= a83[62];
					226:word <= a83[63];
					225:word <= a83[64];
					224:word <= a83[65];
					223:word <= a83[66];
					222:word <= a83[67];
					221:word <= a83[68];
					220:word <= a83[69];
					219:word <= a83[70];
					218:word <= a83[71];
					217:word <= a83[72];
					216:word <= a83[73];
					215:word <= a83[74];
					214:word <= a83[75];
					213:word <= a83[76];
					212:word <= a83[77];
					211:word <= a83[78];
					default:word <= a83[79];
					endcase
				end
				124:begin
				case(x)
					290:word <= a84[0];
					289:word <= a84[1];
					287:word <= a84[2];
					286:word <= a84[3];
					285:word <= a84[4];
					284:word <= a84[5];
					283:word <= a84[6];
					282:word <= a84[7];
					281:word <= a84[8];
					280:word <= a84[9];
					279:word <= a84[10];
					278:word <= a84[11];
					277:word <= a84[12];
					276:word <= a84[13];
					275:word <= a84[14];
					274:word <= a84[15];
					273:word <= a84[16];
					272:word <= a84[17];
					271:word <= a84[18];
					270:word <= a84[19];
					269:word <= a84[20];
					268:word <= a84[21];
					267:word <= a84[22];
					266:word <= a84[23];
					265:word <= a84[24];
					264:word <= a84[25];
					263:word <= a84[26];
					262:word <= a84[27];
					261:word <= a84[28];
					260:word <= a84[29];
					259:word <= a84[30];
					258:word <= a84[31];
					257:word <= a84[32];
					256:word <= a84[33];
					255:word <= a84[34];
					254:word <= a84[35];
					253:word <= a84[36];
					252:word <= a84[37];
					251:word <= a84[38];
					250:word <= a84[39];
					249:word <= a84[40];
					248:word <= a84[41];
					247:word <= a84[42];
					246:word <= a84[43];
					245:word <= a84[44];
					244:word <= a84[45];
					243:word <= a84[46];
					242:word <= a84[47];
					241:word <= a84[48];
					240:word <= a84[49];
					239:word <= a84[50];
					238:word <= a84[51];
					237:word <= a84[52];
					236:word <= a84[53];
					235:word <= a84[54];
					234:word <= a84[55];
					233:word <= a84[56];
					232:word <= a84[57];
					231:word <= a84[58];
					230:word <= a84[59];
					229:word <= a84[60];
					228:word <= a84[61];
					227:word <= a84[62];
					226:word <= a84[63];
					225:word <= a84[64];
					224:word <= a84[65];
					223:word <= a84[66];
					222:word <= a84[67];
					221:word <= a84[68];
					220:word <= a84[69];
					219:word <= a84[70];
					218:word <= a84[71];
					217:word <= a84[72];
					216:word <= a84[73];
					215:word <= a84[74];
					214:word <= a84[75];
					213:word <= a84[76];
					212:word <= a84[77];
					211:word <= a84[78];
					default:word <= a84[79];
					endcase
				end
				125:begin
				case(x)
					290:word <= a85[0];
					289:word <= a85[1];
					287:word <= a85[2];
					286:word <= a85[3];
					285:word <= a85[4];
					284:word <= a85[5];
					283:word <= a85[6];
					282:word <= a85[7];
					281:word <= a85[8];
					280:word <= a85[9];
					279:word <= a85[10];
					278:word <= a85[11];
					277:word <= a85[12];
					276:word <= a85[13];
					275:word <= a85[14];
					274:word <= a85[15];
					273:word <= a85[16];
					272:word <= a85[17];
					271:word <= a85[18];
					270:word <= a85[19];
					269:word <= a85[20];
					268:word <= a85[21];
					267:word <= a85[22];
					266:word <= a85[23];
					265:word <= a85[24];
					264:word <= a85[25];
					263:word <= a85[26];
					262:word <= a85[27];
					261:word <= a85[28];
					260:word <= a85[29];
					259:word <= a85[30];
					258:word <= a85[31];
					257:word <= a85[32];
					256:word <= a85[33];
					255:word <= a85[34];
					254:word <= a85[35];
					253:word <= a85[36];
					252:word <= a85[37];
					251:word <= a85[38];
					250:word <= a85[39];
					249:word <= a85[40];
					248:word <= a85[41];
					247:word <= a85[42];
					246:word <= a85[43];
					245:word <= a85[44];
					244:word <= a85[45];
					243:word <= a85[46];
					242:word <= a85[47];
					241:word <= a85[48];
					240:word <= a85[49];
					239:word <= a85[50];
					238:word <= a85[51];
					237:word <= a85[52];
					236:word <= a85[53];
					235:word <= a85[54];
					234:word <= a85[55];
					233:word <= a85[56];
					232:word <= a85[57];
					231:word <= a85[58];
					230:word <= a85[59];
					229:word <= a85[60];
					228:word <= a85[61];
					227:word <= a85[62];
					226:word <= a85[63];
					225:word <= a85[64];
					224:word <= a85[65];
					223:word <= a85[66];
					222:word <= a85[67];
					221:word <= a85[68];
					220:word <= a85[69];
					219:word <= a85[70];
					218:word <= a85[71];
					217:word <= a85[72];
					216:word <= a85[73];
					215:word <= a85[74];
					214:word <= a85[75];
					213:word <= a85[76];
					212:word <= a85[77];
					211:word <= a85[78];
					default:word <= a85[79];
					endcase
				end
				126:begin
				case(x)
					290:word <= a86[0];
					289:word <= a86[1];
					287:word <= a86[2];
					286:word <= a86[3];
					285:word <= a86[4];
					284:word <= a86[5];
					283:word <= a86[6];
					282:word <= a86[7];
					281:word <= a86[8];
					280:word <= a86[9];
					279:word <= a86[10];
					278:word <= a86[11];
					277:word <= a86[12];
					276:word <= a86[13];
					275:word <= a86[14];
					274:word <= a86[15];
					273:word <= a86[16];
					272:word <= a86[17];
					271:word <= a86[18];
					270:word <= a86[19];
					269:word <= a86[20];
					268:word <= a86[21];
					267:word <= a86[22];
					266:word <= a86[23];
					265:word <= a86[24];
					264:word <= a86[25];
					263:word <= a86[26];
					262:word <= a86[27];
					261:word <= a86[28];
					260:word <= a86[29];
					259:word <= a86[30];
					258:word <= a86[31];
					257:word <= a86[32];
					256:word <= a86[33];
					255:word <= a86[34];
					254:word <= a86[35];
					253:word <= a86[36];
					252:word <= a86[37];
					251:word <= a86[38];
					250:word <= a86[39];
					249:word <= a86[40];
					248:word <= a86[41];
					247:word <= a86[42];
					246:word <= a86[43];
					245:word <= a86[44];
					244:word <= a86[45];
					243:word <= a86[46];
					242:word <= a86[47];
					241:word <= a86[48];
					240:word <= a86[49];
					239:word <= a86[50];
					238:word <= a86[51];
					237:word <= a86[52];
					236:word <= a86[53];
					235:word <= a86[54];
					234:word <= a86[55];
					233:word <= a86[56];
					232:word <= a86[57];
					231:word <= a86[58];
					230:word <= a86[59];
					229:word <= a86[60];
					228:word <= a86[61];
					227:word <= a86[62];
					226:word <= a86[63];
					225:word <= a86[64];
					224:word <= a86[65];
					223:word <= a86[66];
					222:word <= a86[67];
					221:word <= a86[68];
					220:word <= a86[69];
					219:word <= a86[70];
					218:word <= a86[71];
					217:word <= a86[72];
					216:word <= a86[73];
					215:word <= a86[74];
					214:word <= a86[75];
					213:word <= a86[76];
					212:word <= a86[77];
					211:word <= a86[78];
					default:word <= a86[79];
					endcase
				end
				127:begin
				case(x)
					290:word <= a87[0];
					289:word <= a87[1];
					287:word <= a87[2];
					286:word <= a87[3];
					285:word <= a87[4];
					284:word <= a87[5];
					283:word <= a87[6];
					282:word <= a87[7];
					281:word <= a87[8];
					280:word <= a87[9];
					279:word <= a87[10];
					278:word <= a87[11];
					277:word <= a87[12];
					276:word <= a87[13];
					275:word <= a87[14];
					274:word <= a87[15];
					273:word <= a87[16];
					272:word <= a87[17];
					271:word <= a87[18];
					270:word <= a87[19];
					269:word <= a87[20];
					268:word <= a87[21];
					267:word <= a87[22];
					266:word <= a87[23];
					265:word <= a87[24];
					264:word <= a87[25];
					263:word <= a87[26];
					262:word <= a87[27];
					261:word <= a87[28];
					260:word <= a87[29];
					259:word <= a87[30];
					258:word <= a87[31];
					257:word <= a87[32];
					256:word <= a87[33];
					255:word <= a87[34];
					254:word <= a87[35];
					253:word <= a87[36];
					252:word <= a87[37];
					251:word <= a87[38];
					250:word <= a87[39];
					249:word <= a87[40];
					248:word <= a87[41];
					247:word <= a87[42];
					246:word <= a87[43];
					245:word <= a87[44];
					244:word <= a87[45];
					243:word <= a87[46];
					242:word <= a87[47];
					241:word <= a87[48];
					240:word <= a87[49];
					239:word <= a87[50];
					238:word <= a87[51];
					237:word <= a87[52];
					236:word <= a87[53];
					235:word <= a87[54];
					234:word <= a87[55];
					233:word <= a87[56];
					232:word <= a87[57];
					231:word <= a87[58];
					230:word <= a87[59];
					229:word <= a87[60];
					228:word <= a87[61];
					227:word <= a87[62];
					226:word <= a87[63];
					225:word <= a87[64];
					224:word <= a87[65];
					223:word <= a87[66];
					222:word <= a87[67];
					221:word <= a87[68];
					220:word <= a87[69];
					219:word <= a87[70];
					218:word <= a87[71];
					217:word <= a87[72];
					216:word <= a87[73];
					215:word <= a87[74];
					214:word <= a87[75];
					213:word <= a87[76];
					212:word <= a87[77];
					211:word <= a87[78];
					default:word <= a87[79];
					endcase
				end
				128:begin
				case(x)
					290:word <= a88[0];
					289:word <= a88[1];
					287:word <= a88[2];
					286:word <= a88[3];
					285:word <= a88[4];
					284:word <= a88[5];
					283:word <= a88[6];
					282:word <= a88[7];
					281:word <= a88[8];
					280:word <= a88[9];
					279:word <= a88[10];
					278:word <= a88[11];
					277:word <= a88[12];
					276:word <= a88[13];
					275:word <= a88[14];
					274:word <= a88[15];
					273:word <= a88[16];
					272:word <= a88[17];
					271:word <= a88[18];
					270:word <= a88[19];
					269:word <= a88[20];
					268:word <= a88[21];
					267:word <= a88[22];
					266:word <= a88[23];
					265:word <= a88[24];
					264:word <= a88[25];
					263:word <= a88[26];
					262:word <= a88[27];
					261:word <= a88[28];
					260:word <= a88[29];
					259:word <= a88[30];
					258:word <= a88[31];
					257:word <= a88[32];
					256:word <= a88[33];
					255:word <= a88[34];
					254:word <= a88[35];
					253:word <= a88[36];
					252:word <= a88[37];
					251:word <= a88[38];
					250:word <= a88[39];
					249:word <= a88[40];
					248:word <= a88[41];
					247:word <= a88[42];
					246:word <= a88[43];
					245:word <= a88[44];
					244:word <= a88[45];
					243:word <= a88[46];
					242:word <= a88[47];
					241:word <= a88[48];
					240:word <= a88[49];
					239:word <= a88[50];
					238:word <= a88[51];
					237:word <= a88[52];
					236:word <= a88[53];
					235:word <= a88[54];
					234:word <= a88[55];
					233:word <= a88[56];
					232:word <= a88[57];
					231:word <= a88[58];
					230:word <= a88[59];
					229:word <= a88[60];
					228:word <= a88[61];
					227:word <= a88[62];
					226:word <= a88[63];
					225:word <= a88[64];
					224:word <= a88[65];
					223:word <= a88[66];
					222:word <= a88[67];
					221:word <= a88[68];
					220:word <= a88[69];
					219:word <= a88[70];
					218:word <= a88[71];
					217:word <= a88[72];
					216:word <= a88[73];
					215:word <= a88[74];
					214:word <= a88[75];
					213:word <= a88[76];
					212:word <= a88[77];
					211:word <= a88[78];
					default:word <= a88[79];
					endcase
				end
				129:begin
				case(x)
					290:word <= a89[0];
					289:word <= a89[1];
					287:word <= a89[2];
					286:word <= a89[3];
					285:word <= a89[4];
					284:word <= a89[5];
					283:word <= a89[6];
					282:word <= a89[7];
					281:word <= a89[8];
					280:word <= a89[9];
					279:word <= a89[10];
					278:word <= a89[11];
					277:word <= a89[12];
					276:word <= a89[13];
					275:word <= a89[14];
					274:word <= a89[15];
					273:word <= a89[16];
					272:word <= a89[17];
					271:word <= a89[18];
					270:word <= a89[19];
					269:word <= a89[20];
					268:word <= a89[21];
					267:word <= a89[22];
					266:word <= a89[23];
					265:word <= a89[24];
					264:word <= a89[25];
					263:word <= a89[26];
					262:word <= a89[27];
					261:word <= a89[28];
					260:word <= a89[29];
					259:word <= a89[30];
					258:word <= a89[31];
					257:word <= a89[32];
					256:word <= a89[33];
					255:word <= a89[34];
					254:word <= a89[35];
					253:word <= a89[36];
					252:word <= a89[37];
					251:word <= a89[38];
					250:word <= a89[39];
					249:word <= a89[40];
					248:word <= a89[41];
					247:word <= a89[42];
					246:word <= a89[43];
					245:word <= a89[44];
					244:word <= a89[45];
					243:word <= a89[46];
					242:word <= a89[47];
					241:word <= a89[48];
					240:word <= a89[49];
					239:word <= a89[50];
					238:word <= a89[51];
					237:word <= a89[52];
					236:word <= a89[53];
					235:word <= a89[54];
					234:word <= a89[55];
					233:word <= a89[56];
					232:word <= a89[57];
					231:word <= a89[58];
					230:word <= a89[59];
					229:word <= a89[60];
					228:word <= a89[61];
					227:word <= a89[62];
					226:word <= a89[63];
					225:word <= a89[64];
					224:word <= a89[65];
					223:word <= a89[66];
					222:word <= a89[67];
					221:word <= a89[68];
					220:word <= a89[69];
					219:word <= a89[70];
					218:word <= a89[71];
					217:word <= a89[72];
					216:word <= a89[73];
					215:word <= a89[74];
					214:word <= a89[75];
					213:word <= a89[76];
					212:word <= a89[77];
					211:word <= a89[78];
					default:word <= a89[79];
					endcase
				end
				130:begin
				case(x)
					290:word <= a90[0];
					289:word <= a90[1];
					287:word <= a90[2];
					286:word <= a90[3];
					285:word <= a90[4];
					284:word <= a90[5];
					283:word <= a90[6];
					282:word <= a90[7];
					281:word <= a90[8];
					280:word <= a90[9];
					279:word <= a90[10];
					278:word <= a90[11];
					277:word <= a90[12];
					276:word <= a90[13];
					275:word <= a90[14];
					274:word <= a90[15];
					273:word <= a90[16];
					272:word <= a90[17];
					271:word <= a90[18];
					270:word <= a90[19];
					269:word <= a90[20];
					268:word <= a90[21];
					267:word <= a90[22];
					266:word <= a90[23];
					265:word <= a90[24];
					264:word <= a90[25];
					263:word <= a90[26];
					262:word <= a90[27];
					261:word <= a90[28];
					260:word <= a90[29];
					259:word <= a90[30];
					258:word <= a90[31];
					257:word <= a90[32];
					256:word <= a90[33];
					255:word <= a90[34];
					254:word <= a90[35];
					253:word <= a90[36];
					252:word <= a90[37];
					251:word <= a90[38];
					250:word <= a90[39];
					249:word <= a90[40];
					248:word <= a90[41];
					247:word <= a90[42];
					246:word <= a90[43];
					245:word <= a90[44];
					244:word <= a90[45];
					243:word <= a90[46];
					242:word <= a90[47];
					241:word <= a90[48];
					240:word <= a90[49];
					239:word <= a90[50];
					238:word <= a90[51];
					237:word <= a90[52];
					236:word <= a90[53];
					235:word <= a90[54];
					234:word <= a90[55];
					233:word <= a90[56];
					232:word <= a90[57];
					231:word <= a90[58];
					230:word <= a90[59];
					229:word <= a90[60];
					228:word <= a90[61];
					227:word <= a90[62];
					226:word <= a90[63];
					225:word <= a90[64];
					224:word <= a90[65];
					223:word <= a90[66];
					222:word <= a90[67];
					221:word <= a90[68];
					220:word <= a90[69];
					219:word <= a90[70];
					218:word <= a90[71];
					217:word <= a90[72];
					216:word <= a90[73];
					215:word <= a90[74];
					214:word <= a90[75];
					213:word <= a90[76];
					212:word <= a90[77];
					211:word <= a90[78];
					default:word <= a90[79];
					endcase
				end

			131:begin
				case(x)
					290:word <= a91[0];
					289:word <= a91[1];
					287:word <= a91[2];
					286:word <= a91[3];
					285:word <= a91[4];
					284:word <= a91[5];
					283:word <= a91[6];
					282:word <= a91[7];
					281:word <= a91[8];
					280:word <= a91[9];
					279:word <= a91[10];
					278:word <= a91[11];
					277:word <= a91[12];
					276:word <= a91[13];
					275:word <= a91[14];
					274:word <= a91[15];
					273:word <= a91[16];
					272:word <= a91[17];
					271:word <= a91[18];
					270:word <= a91[19];
					269:word <= a91[20];
					268:word <= a91[21];
					267:word <= a91[22];
					266:word <= a91[23];
					265:word <= a91[24];
					264:word <= a91[25];
					263:word <= a91[26];
					262:word <= a91[27];
					261:word <= a91[28];
					260:word <= a91[29];
					259:word <= a91[30];
					258:word <= a91[31];
					257:word <= a91[32];
					256:word <= a91[33];
					255:word <= a91[34];
					254:word <= a91[35];
					253:word <= a91[36];
					252:word <= a91[37];
					251:word <= a91[38];
					250:word <= a91[39];
					249:word <= a91[40];
					248:word <= a91[41];
					247:word <= a91[42];
					246:word <= a91[43];
					245:word <= a91[44];
					244:word <= a91[45];
					243:word <= a91[46];
					242:word <= a91[47];
					241:word <= a91[48];
					240:word <= a91[49];
					239:word <= a91[50];
					238:word <= a91[51];
					237:word <= a91[52];
					236:word <= a91[53];
					235:word <= a91[54];
					234:word <= a91[55];
					233:word <= a91[56];
					232:word <= a91[57];
					231:word <= a91[58];
					230:word <= a91[59];
					229:word <= a91[60];
					228:word <= a91[61];
					227:word <= a91[62];
					226:word <= a91[63];
					225:word <= a91[64];
					224:word <= a91[65];
					223:word <= a91[66];
					222:word <= a91[67];
					221:word <= a91[68];
					220:word <= a91[69];
					219:word <= a91[70];
					218:word <= a91[71];
					217:word <= a91[72];
					216:word <= a91[73];
					215:word <= a91[74];
					214:word <= a91[75];
					213:word <= a91[76];
					212:word <= a91[77];
					211:word <= a91[78];
					default:word <= a91[79];
					endcase
				end
				132:begin
				case(x)
					290:word <= a92[0];
					289:word <= a92[1];
					287:word <= a92[2];
					286:word <= a92[3];
					285:word <= a92[4];
					284:word <= a92[5];
					283:word <= a92[6];
					282:word <= a92[7];
					281:word <= a92[8];
					280:word <= a92[9];
					279:word <= a92[10];
					278:word <= a92[11];
					277:word <= a92[12];
					276:word <= a92[13];
					275:word <= a92[14];
					274:word <= a92[15];
					273:word <= a92[16];
					272:word <= a92[17];
					271:word <= a92[18];
					270:word <= a92[19];
					269:word <= a92[20];
					268:word <= a92[21];
					267:word <= a92[22];
					266:word <= a92[23];
					265:word <= a92[24];
					264:word <= a92[25];
					263:word <= a92[26];
					262:word <= a92[27];
					261:word <= a92[28];
					260:word <= a92[29];
					259:word <= a92[30];
					258:word <= a92[31];
					257:word <= a92[32];
					256:word <= a92[33];
					255:word <= a92[34];
					254:word <= a92[35];
					253:word <= a92[36];
					252:word <= a92[37];
					251:word <= a92[38];
					250:word <= a92[39];
					249:word <= a92[40];
					248:word <= a92[41];
					247:word <= a92[42];
					246:word <= a92[43];
					245:word <= a92[44];
					244:word <= a92[45];
					243:word <= a92[46];
					242:word <= a92[47];
					241:word <= a92[48];
					240:word <= a92[49];
					239:word <= a92[50];
					238:word <= a92[51];
					237:word <= a92[52];
					236:word <= a92[53];
					235:word <= a92[54];
					234:word <= a92[55];
					233:word <= a92[56];
					232:word <= a92[57];
					231:word <= a92[58];
					230:word <= a92[59];
					229:word <= a92[60];
					228:word <= a92[61];
					227:word <= a92[62];
					226:word <= a92[63];
					225:word <= a92[64];
					224:word <= a92[65];
					223:word <= a92[66];
					222:word <= a92[67];
					221:word <= a92[68];
					220:word <= a92[69];
					219:word <= a92[70];
					218:word <= a92[71];
					217:word <= a92[72];
					216:word <= a92[73];
					215:word <= a92[74];
					214:word <= a92[75];
					213:word <= a92[76];
					212:word <= a92[77];
					211:word <= a92[78];
					default:word <= a92[79];
					endcase
				end
				133:begin
				case(x)
					290:word <= a93[0];
					289:word <= a93[1];
					287:word <= a93[2];
					286:word <= a93[3];
					285:word <= a93[4];
					284:word <= a93[5];
					283:word <= a93[6];
					282:word <= a93[7];
					281:word <= a93[8];
					280:word <= a93[9];
					279:word <= a93[10];
					278:word <= a93[11];
					277:word <= a93[12];
					276:word <= a93[13];
					275:word <= a93[14];
					274:word <= a93[15];
					273:word <= a93[16];
					272:word <= a93[17];
					271:word <= a93[18];
					270:word <= a93[19];
					269:word <= a93[20];
					268:word <= a93[21];
					267:word <= a93[22];
					266:word <= a93[23];
					265:word <= a93[24];
					264:word <= a93[25];
					263:word <= a93[26];
					262:word <= a93[27];
					261:word <= a93[28];
					260:word <= a93[29];
					259:word <= a93[30];
					258:word <= a93[31];
					257:word <= a93[32];
					256:word <= a93[33];
					255:word <= a93[34];
					254:word <= a93[35];
					253:word <= a93[36];
					252:word <= a93[37];
					251:word <= a93[38];
					250:word <= a93[39];
					249:word <= a93[40];
					248:word <= a93[41];
					247:word <= a93[42];
					246:word <= a93[43];
					245:word <= a93[44];
					244:word <= a93[45];
					243:word <= a93[46];
					242:word <= a93[47];
					241:word <= a93[48];
					240:word <= a93[49];
					239:word <= a93[50];
					238:word <= a93[51];
					237:word <= a93[52];
					236:word <= a93[53];
					235:word <= a93[54];
					234:word <= a93[55];
					233:word <= a93[56];
					232:word <= a93[57];
					231:word <= a93[58];
					230:word <= a93[59];
					229:word <= a93[60];
					228:word <= a93[61];
					227:word <= a93[62];
					226:word <= a93[63];
					225:word <= a93[64];
					224:word <= a93[65];
					223:word <= a93[66];
					222:word <= a93[67];
					221:word <= a93[68];
					220:word <= a93[69];
					219:word <= a93[70];
					218:word <= a93[71];
					217:word <= a93[72];
					216:word <= a93[73];
					215:word <= a93[74];
					214:word <= a93[75];
					213:word <= a93[76];
					212:word <= a93[77];
					211:word <= a93[78];
					default:word <= a93[79];
					endcase
				end
				134:begin
				case(x)
					290:word <= a94[0];
					289:word <= a94[1];
					287:word <= a94[2];
					286:word <= a94[3];
					285:word <= a94[4];
					284:word <= a94[5];
					283:word <= a94[6];
					282:word <= a94[7];
					281:word <= a94[8];
					280:word <= a94[9];
					279:word <= a94[10];
					278:word <= a94[11];
					277:word <= a94[12];
					276:word <= a94[13];
					275:word <= a94[14];
					274:word <= a94[15];
					273:word <= a94[16];
					272:word <= a94[17];
					271:word <= a94[18];
					270:word <= a94[19];
					269:word <= a94[20];
					268:word <= a94[21];
					267:word <= a94[22];
					266:word <= a94[23];
					265:word <= a94[24];
					264:word <= a94[25];
					263:word <= a94[26];
					262:word <= a94[27];
					261:word <= a94[28];
					260:word <= a94[29];
					259:word <= a94[30];
					258:word <= a94[31];
					257:word <= a94[32];
					256:word <= a94[33];
					255:word <= a94[34];
					254:word <= a94[35];
					253:word <= a94[36];
					252:word <= a94[37];
					251:word <= a94[38];
					250:word <= a94[39];
					249:word <= a94[40];
					248:word <= a94[41];
					247:word <= a94[42];
					246:word <= a94[43];
					245:word <= a94[44];
					244:word <= a94[45];
					243:word <= a94[46];
					242:word <= a94[47];
					241:word <= a94[48];
					240:word <= a94[49];
					239:word <= a94[50];
					238:word <= a94[51];
					237:word <= a94[52];
					236:word <= a94[53];
					235:word <= a94[54];
					234:word <= a94[55];
					233:word <= a94[56];
					232:word <= a94[57];
					231:word <= a94[58];
					230:word <= a94[59];
					229:word <= a94[60];
					228:word <= a94[61];
					227:word <= a94[62];
					226:word <= a94[63];
					225:word <= a94[64];
					224:word <= a94[65];
					223:word <= a94[66];
					222:word <= a94[67];
					221:word <= a94[68];
					220:word <= a94[69];
					219:word <= a94[70];
					218:word <= a94[71];
					217:word <= a94[72];
					216:word <= a94[73];
					215:word <= a94[74];
					214:word <= a94[75];
					213:word <= a94[76];
					212:word <= a94[77];
					211:word <= a94[78];
					default:word <= a94[79];
					endcase
				end
				135:begin
				case(x)
					290:word <= a95[0];
					289:word <= a95[1];
					287:word <= a95[2];
					286:word <= a95[3];
					285:word <= a95[4];
					284:word <= a95[5];
					283:word <= a95[6];
					282:word <= a95[7];
					281:word <= a95[8];
					280:word <= a95[9];
					279:word <= a95[10];
					278:word <= a95[11];
					277:word <= a95[12];
					276:word <= a95[13];
					275:word <= a95[14];
					274:word <= a95[15];
					273:word <= a95[16];
					272:word <= a95[17];
					271:word <= a95[18];
					270:word <= a95[19];
					269:word <= a95[20];
					268:word <= a95[21];
					267:word <= a95[22];
					266:word <= a95[23];
					265:word <= a95[24];
					264:word <= a95[25];
					263:word <= a95[26];
					262:word <= a95[27];
					261:word <= a95[28];
					260:word <= a95[29];
					259:word <= a95[30];
					258:word <= a95[31];
					257:word <= a95[32];
					256:word <= a95[33];
					255:word <= a95[34];
					254:word <= a95[35];
					253:word <= a95[36];
					252:word <= a95[37];
					251:word <= a95[38];
					250:word <= a95[39];
					249:word <= a95[40];
					248:word <= a95[41];
					247:word <= a95[42];
					246:word <= a95[43];
					245:word <= a95[44];
					244:word <= a95[45];
					243:word <= a95[46];
					242:word <= a95[47];
					241:word <= a95[48];
					240:word <= a95[49];
					239:word <= a95[50];
					238:word <= a95[51];
					237:word <= a95[52];
					236:word <= a95[53];
					235:word <= a95[54];
					234:word <= a95[55];
					233:word <= a95[56];
					232:word <= a95[57];
					231:word <= a95[58];
					230:word <= a95[59];
					229:word <= a95[60];
					228:word <= a95[61];
					227:word <= a95[62];
					226:word <= a95[63];
					225:word <= a95[64];
					224:word <= a95[65];
					223:word <= a95[66];
					222:word <= a95[67];
					221:word <= a95[68];
					220:word <= a95[69];
					219:word <= a95[70];
					218:word <= a95[71];
					217:word <= a95[72];
					216:word <= a95[73];
					215:word <= a95[74];
					214:word <= a95[75];
					213:word <= a95[76];
					212:word <= a95[77];
					211:word <= a95[78];
					default:word <= a95[79];
					endcase
				end
				136:begin
				case(x)
					290:word <= a96[0];
					289:word <= a96[1];
					287:word <= a96[2];
					286:word <= a96[3];
					285:word <= a96[4];
					284:word <= a96[5];
					283:word <= a96[6];
					282:word <= a96[7];
					281:word <= a96[8];
					280:word <= a96[9];
					279:word <= a96[10];
					278:word <= a96[11];
					277:word <= a96[12];
					276:word <= a96[13];
					275:word <= a96[14];
					274:word <= a96[15];
					273:word <= a96[16];
					272:word <= a96[17];
					271:word <= a96[18];
					270:word <= a96[19];
					269:word <= a96[20];
					268:word <= a96[21];
					267:word <= a96[22];
					266:word <= a96[23];
					265:word <= a96[24];
					264:word <= a96[25];
					263:word <= a96[26];
					262:word <= a96[27];
					261:word <= a96[28];
					260:word <= a96[29];
					259:word <= a96[30];
					258:word <= a96[31];
					257:word <= a96[32];
					256:word <= a96[33];
					255:word <= a96[34];
					254:word <= a96[35];
					253:word <= a96[36];
					252:word <= a96[37];
					251:word <= a96[38];
					250:word <= a96[39];
					249:word <= a96[40];
					248:word <= a96[41];
					247:word <= a96[42];
					246:word <= a96[43];
					245:word <= a96[44];
					244:word <= a96[45];
					243:word <= a96[46];
					242:word <= a96[47];
					241:word <= a96[48];
					240:word <= a96[49];
					239:word <= a96[50];
					238:word <= a96[51];
					237:word <= a96[52];
					236:word <= a96[53];
					235:word <= a96[54];
					234:word <= a96[55];
					233:word <= a96[56];
					232:word <= a96[57];
					231:word <= a96[58];
					230:word <= a96[59];
					229:word <= a96[60];
					228:word <= a96[61];
					227:word <= a96[62];
					226:word <= a96[63];
					225:word <= a96[64];
					224:word <= a96[65];
					223:word <= a96[66];
					222:word <= a96[67];
					221:word <= a96[68];
					220:word <= a96[69];
					219:word <= a96[70];
					218:word <= a96[71];
					217:word <= a96[72];
					216:word <= a96[73];
					215:word <= a96[74];
					214:word <= a96[75];
					213:word <= a96[76];
					212:word <= a96[77];
					211:word <= a96[78];
					default:word <= a96[79];
					endcase
				end
				137:begin
				case(x)
					290:word <= a97[0];
					289:word <= a97[1];
					287:word <= a97[2];
					286:word <= a97[3];
					285:word <= a97[4];
					284:word <= a97[5];
					283:word <= a97[6];
					282:word <= a97[7];
					281:word <= a97[8];
					280:word <= a97[9];
					279:word <= a97[10];
					278:word <= a97[11];
					277:word <= a97[12];
					276:word <= a97[13];
					275:word <= a97[14];
					274:word <= a97[15];
					273:word <= a97[16];
					272:word <= a97[17];
					271:word <= a97[18];
					270:word <= a97[19];
					269:word <= a97[20];
					268:word <= a97[21];
					267:word <= a97[22];
					266:word <= a97[23];
					265:word <= a97[24];
					264:word <= a97[25];
					263:word <= a97[26];
					262:word <= a97[27];
					261:word <= a97[28];
					260:word <= a97[29];
					259:word <= a97[30];
					258:word <= a97[31];
					257:word <= a97[32];
					256:word <= a97[33];
					255:word <= a97[34];
					254:word <= a97[35];
					253:word <= a97[36];
					252:word <= a97[37];
					251:word <= a97[38];
					250:word <= a97[39];
					249:word <= a97[40];
					248:word <= a97[41];
					247:word <= a97[42];
					246:word <= a97[43];
					245:word <= a97[44];
					244:word <= a97[45];
					243:word <= a97[46];
					242:word <= a97[47];
					241:word <= a97[48];
					240:word <= a97[49];
					239:word <= a97[50];
					238:word <= a97[51];
					237:word <= a97[52];
					236:word <= a97[53];
					235:word <= a97[54];
					234:word <= a97[55];
					233:word <= a97[56];
					232:word <= a97[57];
					231:word <= a97[58];
					230:word <= a97[59];
					229:word <= a97[60];
					228:word <= a97[61];
					227:word <= a97[62];
					226:word <= a97[63];
					225:word <= a97[64];
					224:word <= a97[65];
					223:word <= a97[66];
					222:word <= a97[67];
					221:word <= a97[68];
					220:word <= a97[69];
					219:word <= a97[70];
					218:word <= a97[71];
					217:word <= a97[72];
					216:word <= a97[73];
					215:word <= a97[74];
					214:word <= a97[75];
					213:word <= a97[76];
					212:word <= a97[77];
					211:word <= a97[78];
					default:word <= a97[79];
					endcase
				end
				138:begin
				case(x)
					290:word <= a98[0];
					289:word <= a98[1];
					287:word <= a98[2];
					286:word <= a98[3];
					285:word <= a98[4];
					284:word <= a98[5];
					283:word <= a98[6];
					282:word <= a98[7];
					281:word <= a98[8];
					280:word <= a98[9];
					279:word <= a98[10];
					278:word <= a98[11];
					277:word <= a98[12];
					276:word <= a98[13];
					275:word <= a98[14];
					274:word <= a98[15];
					273:word <= a98[16];
					272:word <= a98[17];
					271:word <= a98[18];
					270:word <= a98[19];
					269:word <= a98[20];
					268:word <= a98[21];
					267:word <= a98[22];
					266:word <= a98[23];
					265:word <= a98[24];
					264:word <= a98[25];
					263:word <= a98[26];
					262:word <= a98[27];
					261:word <= a98[28];
					260:word <= a98[29];
					259:word <= a98[30];
					258:word <= a98[31];
					257:word <= a98[32];
					256:word <= a98[33];
					255:word <= a98[34];
					254:word <= a98[35];
					253:word <= a98[36];
					252:word <= a98[37];
					251:word <= a98[38];
					250:word <= a98[39];
					249:word <= a98[40];
					248:word <= a98[41];
					247:word <= a98[42];
					246:word <= a98[43];
					245:word <= a98[44];
					244:word <= a98[45];
					243:word <= a98[46];
					242:word <= a98[47];
					241:word <= a98[48];
					240:word <= a98[49];
					239:word <= a98[50];
					238:word <= a98[51];
					237:word <= a98[52];
					236:word <= a98[53];
					235:word <= a98[54];
					234:word <= a98[55];
					233:word <= a98[56];
					232:word <= a98[57];
					231:word <= a98[58];
					230:word <= a98[59];
					229:word <= a98[60];
					228:word <= a98[61];
					227:word <= a98[62];
					226:word <= a98[63];
					225:word <= a98[64];
					224:word <= a98[65];
					223:word <= a98[66];
					222:word <= a98[67];
					221:word <= a98[68];
					220:word <= a98[69];
					219:word <= a98[70];
					218:word <= a98[71];
					217:word <= a98[72];
					216:word <= a98[73];
					215:word <= a98[74];
					214:word <= a98[75];
					213:word <= a98[76];
					212:word <= a98[77];
					211:word <= a98[78];
					default:word <= a98[79];
					endcase
				end
				139:begin
				case(x)
					290:word <= a99[0];
					289:word <= a99[1];
					287:word <= a99[2];
					286:word <= a99[3];
					285:word <= a99[4];
					284:word <= a99[5];
					283:word <= a99[6];
					282:word <= a99[7];
					281:word <= a99[8];
					280:word <= a99[9];
					279:word <= a99[10];
					278:word <= a99[11];
					277:word <= a99[12];
					276:word <= a99[13];
					275:word <= a99[14];
					274:word <= a99[15];
					273:word <= a99[16];
					272:word <= a99[17];
					271:word <= a99[18];
					270:word <= a99[19];
					269:word <= a99[20];
					268:word <= a99[21];
					267:word <= a99[22];
					266:word <= a99[23];
					265:word <= a99[24];
					264:word <= a99[25];
					263:word <= a99[26];
					262:word <= a99[27];
					261:word <= a99[28];
					260:word <= a99[29];
					259:word <= a99[30];
					258:word <= a99[31];
					257:word <= a99[32];
					256:word <= a99[33];
					255:word <= a99[34];
					254:word <= a99[35];
					253:word <= a99[36];
					252:word <= a99[37];
					251:word <= a99[38];
					250:word <= a99[39];
					249:word <= a99[40];
					248:word <= a99[41];
					247:word <= a99[42];
					246:word <= a99[43];
					245:word <= a99[44];
					244:word <= a99[45];
					243:word <= a99[46];
					242:word <= a99[47];
					241:word <= a99[48];
					240:word <= a99[49];
					239:word <= a99[50];
					238:word <= a99[51];
					237:word <= a99[52];
					236:word <= a99[53];
					235:word <= a99[54];
					234:word <= a99[55];
					233:word <= a99[56];
					232:word <= a99[57];
					231:word <= a99[58];
					230:word <= a99[59];
					229:word <= a99[60];
					228:word <= a99[61];
					227:word <= a99[62];
					226:word <= a99[63];
					225:word <= a99[64];
					224:word <= a99[65];
					223:word <= a99[66];
					222:word <= a99[67];
					221:word <= a99[68];
					220:word <= a99[69];
					219:word <= a99[70];
					218:word <= a99[71];
					217:word <= a99[72];
					216:word <= a99[73];
					215:word <= a99[74];
					214:word <= a99[75];
					213:word <= a99[76];
					212:word <= a99[77];
					211:word <= a99[78];
					default:word <= a99[79];
					endcase
				end
				140:begin
				case(x)
					290:word <= a100[0];
					289:word <= a100[1];
					287:word <= a100[2];
					286:word <= a100[3];
					285:word <= a100[4];
					284:word <= a100[5];
					283:word <= a100[6];
					282:word <= a100[7];
					281:word <= a100[8];
					280:word <= a100[9];
					279:word <= a100[10];
					278:word <= a100[11];
					277:word <= a100[12];
					276:word <= a100[13];
					275:word <= a100[14];
					274:word <= a100[15];
					273:word <= a100[16];
					272:word <= a100[17];
					271:word <= a100[18];
					270:word <= a100[19];
					269:word <= a100[20];
					268:word <= a100[21];
					267:word <= a100[22];
					266:word <= a100[23];
					265:word <= a100[24];
					264:word <= a100[25];
					263:word <= a100[26];
					262:word <= a100[27];
					261:word <= a100[28];
					260:word <= a100[29];
					259:word <= a100[30];
					258:word <= a100[31];
					257:word <= a100[32];
					256:word <= a100[33];
					255:word <= a100[34];
					254:word <= a100[35];
					253:word <= a100[36];
					252:word <= a100[37];
					251:word <= a100[38];
					250:word <= a100[39];
					249:word <= a100[40];
					248:word <= a100[41];
					247:word <= a100[42];
					246:word <= a100[43];
					245:word <= a100[44];
					244:word <= a100[45];
					243:word <= a100[46];
					242:word <= a100[47];
					241:word <= a100[48];
					240:word <= a100[49];
					239:word <= a100[50];
					238:word <= a100[51];
					237:word <= a100[52];
					236:word <= a100[53];
					235:word <= a100[54];
					234:word <= a100[55];
					233:word <= a100[56];
					232:word <= a100[57];
					231:word <= a100[58];
					230:word <= a100[59];
					229:word <= a100[60];
					228:word <= a100[61];
					227:word <= a100[62];
					226:word <= a100[63];
					225:word <= a100[64];
					224:word <= a100[65];
					223:word <= a100[66];
					222:word <= a100[67];
					221:word <= a100[68];
					220:word <= a100[69];
					219:word <= a100[70];
					218:word <= a100[71];
					217:word <= a100[72];
					216:word <= a100[73];
					215:word <= a100[74];
					214:word <= a100[75];
					213:word <= a100[76];
					212:word <= a100[77];
					211:word <= a100[78];
					default:word <= a100[79];
					endcase
				end
				endcase
			end
end
endmodule
